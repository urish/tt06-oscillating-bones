magic
tech sky130A
magscale 1 2
timestamp 1712764311
<< metal1 >>
rect -747 12037 379 12147
rect -4413 11757 -3185 11867
rect -747 11851 -637 12037
rect 1686 12001 3349 12111
rect -4413 10551 -4303 11757
rect -1880 11741 -637 11851
rect 3239 11311 3349 12001
rect 3239 11201 3869 11311
rect 5174 11205 6075 11315
rect -7446 10426 -6488 10526
rect -5208 10441 -4303 10551
rect -7446 8304 -7346 10426
rect 5965 9505 6075 11205
rect 5965 9395 6953 9505
rect 8270 9421 8665 9531
rect -9912 8198 -9286 8298
rect -7966 8204 -7346 8304
rect -9912 5348 -9812 8198
rect 8555 6919 8665 9421
rect 8555 6809 9381 6919
rect 10704 6783 11057 6893
rect 10947 5549 11057 6783
rect 10947 5439 12569 5549
rect -12608 5238 -11300 5338
rect -10042 5248 -9812 5348
rect -12608 1916 -12508 5238
rect 12459 3701 12569 5439
rect 10736 3576 10930 3676
rect 12285 3591 12569 3701
rect -12608 1816 -12382 1916
rect -11064 1836 -10728 1936
rect -10828 -1648 -10728 1836
rect 10736 128 10836 3576
rect 10736 28 11510 128
rect 12804 38 13060 138
rect -12640 -1750 -12354 -1650
rect -11032 -1748 -10728 -1648
rect -12640 -5080 -12540 -1750
rect 12960 -3388 13060 38
rect -12640 -5180 -11342 -5080
rect -10010 -5164 -9712 -5064
rect -9812 -8028 -9712 -5164
rect 8706 -6706 9392 -6606
rect 10852 -6612 10952 -3410
rect 12266 -3488 13060 -3388
rect -9812 -8128 -9298 -8028
rect -7996 -8118 -7292 -8018
rect -7392 -10254 -7292 -8118
rect 8706 -9244 8806 -6706
rect 10714 -6712 10952 -6612
rect 5744 -9354 6964 -9254
rect 8280 -9344 8806 -9244
rect -7392 -10354 -6550 -10254
rect -5200 -10334 -4740 -10234
rect -4840 -11540 -4740 -10334
rect 2354 -11118 3856 -11018
rect 5744 -11034 5844 -9354
rect -4840 -11640 -3194 -11540
rect -1870 -11658 -708 -11558
rect -808 -11830 -708 -11658
rect -808 -11930 376 -11830
rect 2354 -11834 2454 -11118
rect 5184 -11134 5844 -11034
rect 1696 -11934 2454 -11834
<< metal2 >>
rect -198 14598 200 14600
rect -380 14594 380 14598
rect -560 14588 560 14594
rect -742 14580 742 14588
rect -922 14570 922 14580
rect -1104 14558 1104 14570
rect -1284 14544 1284 14558
rect -1464 14526 1464 14544
rect -1644 14508 1644 14526
rect -1824 14486 1824 14508
rect -2004 14462 2004 14486
rect -2184 14436 2184 14462
rect -2362 14408 2362 14436
rect -2540 14376 2540 14408
rect -2720 14344 2720 14376
rect -2898 14308 2898 14344
rect -3074 14272 3074 14308
rect -3252 14232 3252 14272
rect -3428 14198 3428 14232
rect -3428 14194 -160 14198
rect 160 14194 3428 14198
rect -3428 14190 -342 14194
rect -3604 14188 -342 14190
rect 342 14190 3428 14194
rect 342 14188 3604 14190
rect -3604 14180 -522 14188
rect -3604 14170 -704 14180
rect -3604 14158 -884 14170
rect -3604 14146 -1064 14158
rect -3780 14144 -1064 14146
rect -3780 14126 -1244 14144
rect -3780 14108 -1424 14126
rect -3780 14100 -1604 14108
rect -3956 14086 -1604 14100
rect -3956 14062 -1784 14086
rect -3956 14052 -1962 14062
rect -4130 14036 -1962 14052
rect -4130 14008 -2140 14036
rect -4130 14002 -2320 14008
rect -4304 13976 -2320 14002
rect -4304 13950 -2498 13976
rect -4476 13944 -2498 13950
rect -4476 13908 -2674 13944
rect -4476 13894 -2852 13908
rect -4648 13872 -2852 13894
rect -4648 13838 -3028 13872
rect -4820 13832 -3028 13838
rect -4820 13790 -3204 13832
rect -4820 13778 -3380 13790
rect -4992 13746 -3380 13778
rect -4992 13716 -3556 13746
rect -5162 13700 -3556 13716
rect -5162 13654 -3730 13700
rect -5332 13652 -3730 13654
rect -5332 13602 -3904 13652
rect -5332 13588 -4076 13602
rect -5500 13550 -4076 13588
rect -5500 13520 -4248 13550
rect -5668 13494 -4248 13520
rect -5668 13450 -4420 13494
rect -5834 13438 -4420 13450
rect -5834 13378 -4592 13438
rect -6000 13316 -4762 13378
rect -6000 13304 -4932 13316
rect -6166 13254 -4932 13304
rect -6166 13228 -5100 13254
rect -6330 13188 -5100 13228
rect -6330 13150 -5268 13188
rect -6494 13120 -5268 13150
rect -6494 13070 -5434 13120
rect -6656 13050 -5434 13070
rect -6656 12988 -5600 13050
rect -3170 12998 -3090 13832
rect 396 13266 476 14188
rect 522 14180 3604 14188
rect 704 14170 3604 14180
rect 884 14158 3604 14170
rect 1064 14146 3604 14158
rect 1064 14144 3780 14146
rect 1244 14126 3780 14144
rect 1424 14108 3780 14126
rect 1604 14100 3780 14108
rect 1604 14086 3956 14100
rect 1784 14062 3956 14086
rect 1962 14052 3956 14062
rect 1962 14036 4130 14052
rect 2140 14008 4130 14036
rect 2320 14002 4130 14008
rect 2320 13976 4304 14002
rect 2498 13950 4304 13976
rect 2498 13944 4476 13950
rect 2674 13908 4476 13944
rect 2852 13894 4476 13908
rect 2852 13872 4648 13894
rect 3028 13838 4648 13872
rect 3028 13832 4820 13838
rect 3204 13790 4820 13832
rect 3380 13778 4820 13790
rect 3380 13746 4992 13778
rect 3556 13716 4992 13746
rect 3556 13700 5162 13716
rect 3730 13654 5162 13700
rect 3730 13652 5332 13654
rect 3884 13602 5332 13652
rect -6816 12978 -5600 12988
rect -6816 12904 -5766 12978
rect -6978 12828 -5930 12904
rect -6978 12818 -6094 12828
rect -7136 12750 -6094 12818
rect -7136 12730 -6256 12750
rect -7294 12670 -6256 12730
rect -7294 12640 -6416 12670
rect -7452 12588 -6416 12640
rect -7452 12548 -6578 12588
rect -7606 12504 -6578 12548
rect -7606 12454 -6736 12504
rect -7762 12418 -6736 12454
rect -7762 12358 -6894 12418
rect -7914 12330 -6894 12358
rect -7914 12260 -7052 12330
rect -8068 12240 -7052 12260
rect -8068 12160 -7206 12240
rect -8218 12148 -7206 12160
rect -8218 12058 -7362 12148
rect -8368 12054 -7362 12058
rect -8368 11958 -7514 12054
rect -8368 11954 -7668 11958
rect -8516 11860 -7668 11954
rect -8516 11848 -7818 11860
rect -8664 11760 -7818 11848
rect -8664 11742 -7968 11760
rect -8808 11658 -7968 11742
rect -6498 11692 -6418 12588
rect 3884 12470 3964 13602
rect 4076 13588 5332 13602
rect 4076 13550 5500 13588
rect 4248 13520 5500 13550
rect 4248 13494 5668 13520
rect 4420 13450 5668 13494
rect 4420 13438 5834 13450
rect 4592 13378 5834 13438
rect 4762 13316 6000 13378
rect 4932 13304 6000 13316
rect 4932 13254 6166 13304
rect 5100 13228 6166 13254
rect 5100 13188 6330 13228
rect 5268 13150 6330 13188
rect 5268 13120 6494 13150
rect 5434 13070 6494 13120
rect 5434 13050 6656 13070
rect 5600 12988 6656 13050
rect 5600 12978 6816 12988
rect 5766 12904 6816 12978
rect 5930 12828 6978 12904
rect 6094 12818 6978 12828
rect 6094 12750 7136 12818
rect 6256 12730 7136 12750
rect 6256 12670 7294 12730
rect 6416 12640 7294 12670
rect 6416 12588 7452 12640
rect 6578 12548 7452 12588
rect 6578 12504 7606 12548
rect 6736 12454 7606 12504
rect 6736 12418 7762 12454
rect 6894 12358 7762 12418
rect 6894 12330 7914 12358
rect 6980 12260 7914 12330
rect 6980 12240 8068 12260
rect -8808 11632 -8116 11658
rect -8954 11554 -8116 11632
rect -8954 11522 -8264 11554
rect -9096 11448 -8264 11522
rect -9096 11408 -8408 11448
rect -9238 11342 -8408 11408
rect -9238 11294 -8554 11342
rect -9378 11232 -8554 11294
rect -9378 11178 -8696 11232
rect -9516 11122 -8696 11178
rect -9516 11060 -8838 11122
rect -9654 11008 -8838 11060
rect -9654 10940 -8978 11008
rect -9790 10894 -8978 10940
rect -9790 10820 -9116 10894
rect -9924 10778 -9116 10820
rect -9924 10696 -9216 10778
rect -10056 10660 -9216 10696
rect -10056 10572 -9390 10660
rect -10188 10540 -9390 10572
rect -10188 10446 -9524 10540
rect -10318 10420 -9524 10446
rect -10318 10318 -9656 10420
rect -10446 10296 -9656 10318
rect -10446 10188 -9788 10296
rect -10572 10172 -9788 10188
rect -10572 10056 -9918 10172
rect -10696 10046 -9918 10056
rect -10696 9924 -10046 10046
rect -10820 9918 -10046 9924
rect -10820 9790 -10172 9918
rect -10940 9788 -10172 9790
rect -10940 9656 -10296 9788
rect -10940 9654 -10420 9656
rect -11060 9524 -10420 9654
rect -11060 9516 -10540 9524
rect -11178 9390 -10540 9516
rect -9296 9462 -9216 10660
rect 292 10726 496 10826
rect -3232 10458 -3070 10558
rect -3232 9520 -3132 10458
rect -198 9998 200 10000
rect 292 9998 392 10726
rect 6980 10680 7060 12240
rect 7206 12160 8068 12240
rect 7206 12148 8218 12160
rect 7362 12058 8218 12148
rect 7362 12054 8368 12058
rect 7514 11958 8368 12054
rect 7668 11954 8368 11958
rect 7668 11860 8516 11954
rect 7818 11848 8516 11860
rect 7818 11760 8664 11848
rect 7968 11742 8664 11760
rect 7968 11658 8808 11742
rect 8116 11632 8808 11658
rect 8116 11554 8954 11632
rect 8264 11522 8954 11554
rect 8264 11448 9096 11522
rect 8408 11408 9096 11448
rect 8408 11342 9238 11408
rect 8554 11294 9238 11342
rect 8554 11232 9378 11294
rect 8696 11178 9378 11232
rect 8696 11122 9516 11178
rect 8838 11060 9516 11122
rect 8838 11008 9654 11060
rect 8978 10940 9654 11008
rect 8978 10894 9790 10940
rect 9116 10820 9790 10894
rect 9116 10778 9924 10820
rect 9254 10696 9924 10778
rect 9254 10660 10056 10696
rect 9390 10572 10056 10660
rect 9390 10540 10188 10572
rect 9524 10446 10188 10540
rect 9524 10420 10318 10446
rect 9656 10318 10318 10420
rect 9656 10296 10446 10318
rect 9788 10188 10446 10296
rect 9788 10172 10572 10188
rect 9918 10056 10572 10172
rect 9918 10046 10696 10056
rect -370 9994 392 9998
rect -542 9986 542 9994
rect -712 9976 712 9986
rect -882 9962 882 9976
rect -1054 9946 1054 9962
rect -1224 9926 1224 9946
rect -1394 9904 1394 9926
rect -1562 9878 1562 9904
rect -1732 9850 1732 9878
rect -1900 9818 1900 9850
rect -2068 9784 2068 9818
rect -2236 9748 2236 9784
rect -2404 9708 2404 9748
rect -2570 9666 2570 9708
rect -2736 9620 2736 9666
rect 3884 9642 3984 10030
rect 10046 9924 10696 10046
rect 10046 9918 10820 9924
rect 10172 9790 10820 9918
rect 10172 9788 10940 9790
rect 10296 9656 10940 9788
rect 10420 9654 10940 9656
rect -2900 9598 2900 9620
rect -2900 9594 -142 9598
rect 142 9594 2900 9598
rect -2900 9586 -312 9594
rect 312 9586 2900 9594
rect -2900 9576 -482 9586
rect 482 9576 2900 9586
rect -2900 9570 -654 9576
rect -3064 9562 -654 9570
rect 654 9570 2900 9576
rect 654 9562 3064 9570
rect -3064 9546 -824 9562
rect 824 9546 3064 9562
rect -3064 9526 -994 9546
rect 994 9526 3064 9546
rect 3884 9542 4052 9642
rect -3064 9520 -1162 9526
rect -3232 9504 -1162 9520
rect 1162 9520 3064 9526
rect 1162 9504 3228 9520
rect -3232 9478 -1332 9504
rect 1332 9478 3228 9504
rect -3232 9466 -1500 9478
rect -3390 9450 -1500 9466
rect 1500 9466 3228 9478
rect 1500 9450 3390 9466
rect -3390 9418 -1668 9450
rect 1668 9418 3390 9450
rect -3390 9408 -1836 9418
rect -11178 9378 -10660 9390
rect -11294 9254 -10660 9378
rect -3550 9384 -1836 9408
rect 1836 9408 3390 9418
rect 1836 9384 3550 9408
rect -3550 9348 -2004 9384
rect 2004 9348 3550 9384
rect -3712 9308 -2170 9348
rect 2170 9308 3712 9348
rect -3712 9286 -2336 9308
rect -3870 9266 -2336 9286
rect 2336 9286 3712 9308
rect 2336 9266 3870 9286
rect -11294 9238 -10778 9254
rect -11408 9116 -10778 9238
rect -11408 9096 -10894 9116
rect -11522 8978 -10894 9096
rect -11522 8954 -11008 8978
rect -11632 8838 -11008 8954
rect -11632 8808 -11122 8838
rect -11742 8696 -11122 8808
rect -11742 8664 -11232 8696
rect -11848 8554 -11232 8664
rect -11848 8516 -11342 8554
rect -11954 8408 -11342 8516
rect -11954 8368 -11448 8408
rect -12058 8264 -11448 8368
rect -12058 8218 -11554 8264
rect -12160 8116 -11554 8218
rect -12160 8068 -11658 8116
rect -12260 7968 -11658 8068
rect -12260 7914 -11760 7968
rect -12358 7818 -11760 7914
rect -12358 7762 -11860 7818
rect -12454 7668 -11860 7762
rect -6498 7706 -6398 9252
rect -3870 9220 -2500 9266
rect 2500 9220 3870 9266
rect 3952 9220 4052 9542
rect 10420 9524 11060 9654
rect 10540 9516 11060 9524
rect 10540 9390 11178 9516
rect 10660 9378 11178 9390
rect 10660 9254 11294 9378
rect -4028 9170 -2664 9220
rect 2664 9170 4052 9220
rect 10778 9238 11294 9254
rect 10778 9174 11408 9238
rect -4028 9152 -2828 9170
rect -4186 9120 -2828 9152
rect 2828 9152 4052 9170
rect 2828 9120 4186 9152
rect -4186 9080 -2990 9120
rect -4340 9066 -2990 9080
rect 2990 9080 4186 9120
rect 9414 9096 11408 9174
rect 9414 9094 11522 9096
rect 2990 9066 4340 9080
rect -4340 9008 -3150 9066
rect 3150 9008 4340 9066
rect -4496 8948 -3312 9008
rect 3312 8948 4496 9008
rect -4496 8930 -3470 8948
rect -4648 8886 -3470 8930
rect 3470 8930 4496 8948
rect 3470 8886 4648 8930
rect -4648 8852 -3628 8886
rect -4800 8820 -3628 8852
rect 3628 8852 4648 8886
rect 3628 8820 4800 8852
rect -4800 8770 -3786 8820
rect -4950 8752 -3786 8770
rect 3786 8770 4800 8820
rect 3786 8752 4950 8770
rect -4950 8686 -3940 8752
rect -5098 8680 -3940 8686
rect 3940 8686 4950 8752
rect 3940 8680 5100 8686
rect -5098 8608 -4096 8680
rect 4096 8608 5100 8680
rect -5098 8600 -4248 8608
rect -5246 8530 -4248 8600
rect 4248 8600 5100 8608
rect 4248 8530 5246 8600
rect -5246 8510 -4400 8530
rect -5392 8452 -4400 8510
rect 4400 8510 5246 8530
rect 4400 8452 5392 8510
rect -5392 8418 -4550 8452
rect -5536 8370 -4550 8418
rect 4550 8418 5392 8452
rect 4550 8370 5536 8418
rect -5536 8324 -4698 8370
rect -5680 8286 -4698 8324
rect 4700 8324 5536 8370
rect 4700 8286 5680 8324
rect -5680 8226 -4846 8286
rect -5820 8200 -4846 8226
rect 4846 8226 5680 8286
rect 4846 8200 5820 8226
rect -5820 8128 -4992 8200
rect -5960 8110 -4992 8128
rect 4992 8128 5820 8200
rect 4992 8110 5960 8128
rect -5960 8026 -5136 8110
rect -6096 8018 -5136 8026
rect 5136 8026 5960 8110
rect 5136 8018 6096 8026
rect -6096 7924 -5280 8018
rect 5280 7924 6096 8018
rect -6096 7922 -5420 7924
rect -6232 7826 -5420 7922
rect 5420 7922 6096 7924
rect 5420 7826 6232 7922
rect -6232 7816 -5560 7826
rect -6366 7728 -5560 7816
rect 5560 7816 6232 7826
rect 5560 7728 6366 7816
rect -6366 7706 -5696 7728
rect -12454 7606 -11958 7668
rect -12548 7514 -11958 7606
rect -6498 7626 -5696 7706
rect 5696 7706 6366 7728
rect 5696 7626 6498 7706
rect -6498 7596 -5832 7626
rect -6628 7522 -5832 7596
rect 5832 7596 6498 7626
rect 5832 7522 6628 7596
rect -12548 7452 -12054 7514
rect -6628 7482 -5966 7522
rect -12640 7362 -12054 7452
rect -6756 7416 -5966 7482
rect 5966 7482 6628 7522
rect 5966 7416 6756 7482
rect -6756 7366 -6098 7416
rect -12640 7294 -12148 7362
rect -12730 7206 -12148 7294
rect -6882 7306 -6098 7366
rect 6098 7366 6756 7416
rect 6098 7306 6882 7366
rect -6882 7248 -6228 7306
rect -12730 7136 -12240 7206
rect -12818 7052 -12240 7136
rect -7006 7196 -6228 7248
rect 6228 7248 6882 7306
rect 6980 7248 7080 8240
rect 9414 8058 9494 9094
rect 10894 8978 11522 9094
rect 11008 8954 11522 8978
rect 11008 8838 11632 8954
rect 11122 8808 11632 8838
rect 11122 8696 11742 8808
rect 11232 8664 11742 8696
rect 11232 8554 11848 8664
rect 11342 8516 11848 8554
rect 11342 8408 11954 8516
rect 11448 8368 11954 8408
rect 11448 8264 12058 8368
rect 11554 8218 12058 8264
rect 11554 8116 12160 8218
rect 11658 8068 12160 8116
rect 11658 7968 12260 8068
rect 11760 7914 12260 7968
rect 11760 7818 12358 7914
rect 11860 7762 12358 7818
rect 11860 7668 12454 7762
rect 11958 7606 12454 7668
rect 11958 7514 12548 7606
rect 12054 7452 12548 7514
rect 12054 7362 12640 7452
rect 6228 7196 7080 7248
rect 12148 7294 12640 7362
rect 12148 7206 12730 7294
rect -7006 7128 -6356 7196
rect -7128 7082 -6356 7128
rect 6356 7128 7080 7196
rect 12240 7136 12730 7206
rect 6356 7082 7128 7128
rect -12818 6978 -12330 7052
rect -12904 6894 -12330 6978
rect -12904 6816 -12418 6894
rect -12988 6736 -12418 6816
rect -12988 6656 -12504 6736
rect -13070 6586 -12504 6656
rect -13070 6506 -11230 6586
rect -13070 6494 -12588 6506
rect -13150 6416 -12588 6494
rect -13150 6330 -12670 6416
rect -13228 6256 -12670 6330
rect -13228 6166 -12750 6256
rect -13304 6094 -12750 6166
rect -9296 6128 -9196 7022
rect -7128 7006 -6482 7082
rect -7248 6966 -6482 7006
rect 6482 7006 7128 7082
rect 12240 7052 12818 7136
rect 6482 6966 7248 7006
rect -7248 6882 -6606 6966
rect -7366 6848 -6606 6882
rect 6606 6882 7248 6966
rect 12330 6978 12818 7052
rect 12330 6894 12904 6978
rect 6606 6848 7366 6882
rect -7366 6756 -6728 6848
rect -7482 6728 -6728 6756
rect 6728 6756 7366 6848
rect 12418 6816 12904 6894
rect 6728 6728 7482 6756
rect 12418 6736 12988 6816
rect -7482 6628 -6848 6728
rect -7596 6606 -6848 6628
rect 6848 6628 7482 6728
rect 12504 6656 12988 6736
rect 6848 6606 7596 6628
rect -7596 6498 -6966 6606
rect -7706 6482 -6966 6498
rect 6966 6498 7596 6606
rect 12504 6578 13070 6656
rect 6966 6482 7706 6498
rect -7706 6366 -7082 6482
rect -7816 6356 -7082 6366
rect 7082 6366 7706 6482
rect 12588 6494 13070 6578
rect 12588 6416 13150 6494
rect 7082 6356 7816 6366
rect -7816 6232 -7196 6356
rect -7922 6228 -7196 6232
rect 7196 6232 7816 6356
rect 12670 6330 13150 6416
rect 12670 6256 13228 6330
rect 7196 6228 7922 6232
rect -7922 6128 -7306 6228
rect -9296 6098 -7306 6128
rect 7306 6098 7922 6228
rect -13304 6000 -12828 6094
rect -9296 6028 -7416 6098
rect -13378 5930 -12828 6000
rect -8026 5966 -7416 6028
rect 7416 6096 7922 6098
rect 12750 6166 13228 6256
rect 7416 5966 8026 6096
rect 12750 6094 13304 6166
rect -8026 5960 -7522 5966
rect -13378 5834 -12904 5930
rect -13450 5766 -12904 5834
rect -8128 5832 -7522 5960
rect 7522 5960 8026 5966
rect 12828 6000 13304 6094
rect 7522 5832 8128 5960
rect 12828 5930 13378 6000
rect -8128 5820 -7626 5832
rect -13450 5668 -12978 5766
rect -8226 5696 -7626 5820
rect 7626 5820 8128 5832
rect 12904 5834 13378 5930
rect 7626 5696 8226 5820
rect 12904 5766 13450 5834
rect -8226 5680 -7728 5696
rect -13520 5600 -12978 5668
rect -13520 5500 -13050 5600
rect -8324 5560 -7728 5680
rect 7728 5680 8226 5696
rect 7728 5618 8324 5680
rect 12978 5668 13450 5766
rect 7728 5560 9514 5618
rect 12978 5600 13520 5668
rect -8324 5536 -7826 5560
rect -13588 5434 -13050 5500
rect -13588 5332 -13120 5434
rect -8418 5420 -7826 5536
rect 7826 5518 9514 5560
rect 7826 5420 8418 5518
rect 13050 5500 13520 5600
rect 13050 5434 13588 5500
rect -8418 5392 -7924 5420
rect -13654 5268 -13120 5332
rect -8510 5280 -7924 5392
rect 7924 5392 8418 5420
rect 7924 5280 8510 5392
rect -13654 5162 -13188 5268
rect -8510 5246 -8018 5280
rect -13716 5100 -13188 5162
rect -8600 5136 -8018 5246
rect 8018 5246 8510 5280
rect 13120 5332 13588 5434
rect 13120 5268 13654 5332
rect 8018 5136 8600 5246
rect -13716 4992 -13254 5100
rect -8600 5098 -8110 5136
rect -13778 4932 -13254 4992
rect -8686 4992 -8110 5098
rect 8110 5098 8600 5136
rect 13188 5162 13654 5268
rect 13188 5100 13716 5162
rect 8110 4992 8686 5098
rect 13254 5020 13716 5100
rect -8686 4950 -8200 4992
rect -13778 4820 -13316 4932
rect -13838 4762 -13316 4820
rect -8770 4846 -8200 4950
rect 8200 4950 8686 4992
rect 12196 4992 13716 5020
rect 8200 4846 8770 4950
rect -8770 4800 -8286 4846
rect -13838 4648 -13378 4762
rect -8852 4698 -8286 4800
rect 8286 4800 8770 4846
rect 12196 4940 13778 4992
rect 12196 4836 12276 4940
rect 13254 4932 13778 4940
rect 13316 4820 13778 4932
rect 8286 4698 8852 4800
rect 13316 4762 13838 4820
rect -8852 4648 -8370 4698
rect -13894 4592 -13378 4648
rect -13894 4476 -13438 4592
rect -8930 4550 -8370 4648
rect 8370 4648 8852 4698
rect 13378 4648 13838 4762
rect 8370 4550 8930 4648
rect 13378 4592 13894 4648
rect -8930 4496 -8452 4550
rect -13950 4420 -13438 4476
rect -13950 4304 -13494 4420
rect -9008 4400 -8452 4496
rect 8452 4496 8930 4550
rect 8452 4400 9008 4496
rect 13438 4476 13894 4592
rect 13438 4420 13950 4476
rect -9008 4340 -8530 4400
rect -14002 4248 -13494 4304
rect -9080 4248 -8530 4340
rect 8530 4340 9008 4400
rect 8530 4248 9080 4340
rect 13494 4304 13950 4420
rect 13494 4248 14002 4304
rect -14002 4130 -13550 4248
rect -9080 4186 -8608 4248
rect -14052 4076 -13550 4130
rect -9152 4096 -8608 4186
rect 8608 4186 9080 4248
rect 8608 4096 9152 4186
rect -14052 3956 -13602 4076
rect -14100 3904 -13602 3956
rect -14100 3780 -13652 3904
rect -14146 3730 -13652 3780
rect -11310 3858 -11210 4066
rect -9152 4028 -8680 4096
rect -9220 3940 -8680 4028
rect 8680 4028 9152 4096
rect 13550 4130 14002 4248
rect 13550 4076 14052 4130
rect 8680 3940 9220 4028
rect -9220 3870 -8752 3940
rect -9286 3858 -8752 3870
rect -11310 3786 -8752 3858
rect 8752 3870 9220 3940
rect 13602 3956 14052 4076
rect 13602 3904 14100 3956
rect 8752 3786 9286 3870
rect -11310 3758 -8820 3786
rect -14146 3604 -13700 3730
rect -9286 3712 -8820 3758
rect -14190 3556 -13700 3604
rect -9348 3628 -8820 3712
rect 8820 3712 9286 3786
rect 13652 3780 14100 3904
rect 13652 3730 14146 3780
rect 8820 3628 9348 3712
rect -14190 3428 -13746 3556
rect -9348 3550 -8886 3628
rect -14232 3380 -13746 3428
rect -9408 3470 -8886 3550
rect 8886 3550 9348 3628
rect 13700 3604 14146 3730
rect 13700 3556 14190 3604
rect 8886 3470 9408 3550
rect -9408 3390 -8948 3470
rect -14232 3352 -13790 3380
rect -14232 3272 -11054 3352
rect -14232 3252 -13790 3272
rect -14272 3204 -13790 3252
rect -14272 3074 -13832 3204
rect -11134 3088 -11054 3272
rect -9466 3312 -8948 3390
rect 8948 3390 9408 3470
rect 13746 3428 14190 3556
rect 8948 3312 9466 3390
rect 13746 3380 14232 3428
rect -9466 3228 -9008 3312
rect -9520 3150 -9008 3228
rect 9008 3228 9466 3312
rect 13790 3252 14232 3380
rect 9008 3150 9520 3228
rect 13790 3204 14272 3252
rect -14308 3028 -13832 3074
rect -9520 3064 -9066 3150
rect -14308 2898 -13872 3028
rect -9570 2990 -9066 3064
rect 9066 3064 9520 3150
rect 13832 3074 14272 3204
rect 9066 2990 9570 3064
rect 13832 3028 14308 3074
rect -9570 2900 -9120 2990
rect -14344 2852 -13872 2898
rect -14344 2720 -13908 2852
rect -9620 2828 -9120 2900
rect 9120 2900 9570 2990
rect 9120 2828 9620 2900
rect 13872 2898 14308 3028
rect 13872 2852 14344 2898
rect -9620 2736 -9170 2828
rect -14376 2674 -13908 2720
rect -14376 2540 -13944 2674
rect -9666 2664 -9170 2736
rect 9170 2736 9620 2828
rect 9170 2664 9666 2736
rect 13908 2720 14344 2852
rect 13908 2674 14376 2720
rect -9666 2570 -9220 2664
rect -14408 2498 -13944 2540
rect -9708 2500 -9220 2570
rect 9220 2570 9666 2664
rect 9220 2500 9708 2570
rect -14408 2362 -13976 2498
rect -9708 2404 -9266 2500
rect -14436 2320 -13976 2362
rect -9748 2336 -9266 2404
rect 9266 2404 9708 2500
rect 13944 2540 14376 2674
rect 13944 2498 14408 2540
rect 9266 2336 9748 2404
rect -14436 2184 -14008 2320
rect -9748 2236 -9308 2336
rect -14462 2140 -14008 2184
rect -9784 2170 -9308 2236
rect 9308 2236 9748 2336
rect 13976 2362 14408 2498
rect 13976 2320 14436 2362
rect 9308 2170 9784 2236
rect -14462 2004 -14036 2140
rect -9784 2068 -9348 2170
rect -14486 1962 -14036 2004
rect -9818 2004 -9348 2068
rect 9348 2068 9784 2170
rect 14008 2184 14436 2320
rect 14008 2140 14462 2184
rect 9348 2004 9818 2068
rect -14486 1824 -14062 1962
rect -9818 1900 -9384 2004
rect -14508 1784 -14062 1824
rect -9850 1836 -9384 1900
rect 9384 1900 9818 2004
rect 14036 2004 14462 2140
rect 14036 1962 14486 2004
rect 9384 1836 9850 1900
rect -14508 1644 -14086 1784
rect -9850 1732 -9418 1836
rect -14526 1604 -14086 1644
rect -9878 1668 -9418 1732
rect 9418 1732 9850 1836
rect 14062 1824 14486 1962
rect 14062 1784 14508 1824
rect 9418 1668 9878 1732
rect -14526 1464 -14108 1604
rect -9878 1562 -9450 1668
rect -14544 1424 -14108 1464
rect -9904 1500 -9450 1562
rect 9450 1562 9878 1668
rect 14086 1644 14508 1784
rect 14086 1604 14526 1644
rect 9450 1500 9904 1562
rect 14108 1556 14526 1604
rect -14544 1284 -14126 1424
rect -9904 1394 -9478 1500
rect -14558 1244 -14126 1284
rect -9926 1332 -9478 1394
rect 9478 1394 9904 1500
rect 11500 1476 14526 1556
rect 9478 1332 9926 1394
rect -14558 1104 -14144 1244
rect -9926 1224 -9504 1332
rect -14570 1064 -14144 1104
rect -9946 1162 -9504 1224
rect 9504 1224 9926 1332
rect 11500 1300 11580 1476
rect 14108 1464 14526 1476
rect 14108 1424 14544 1464
rect 14126 1284 14544 1424
rect 14126 1244 14558 1284
rect 9504 1162 9946 1224
rect -14570 922 -14158 1064
rect -9946 1054 -9526 1162
rect -14580 884 -14158 922
rect -9962 994 -9526 1054
rect 9526 1054 9946 1162
rect 14144 1104 14558 1244
rect 14144 1064 14570 1104
rect 9526 994 9962 1054
rect -14580 742 -14170 884
rect -9962 882 -9546 994
rect -14588 704 -14170 742
rect -9976 824 -9546 882
rect 9546 882 9962 994
rect 14158 922 14570 1064
rect 14158 884 14580 922
rect 9546 824 9976 882
rect -9976 712 -9562 824
rect -14588 560 -14180 704
rect -9986 654 -9562 712
rect 9562 712 9976 824
rect 14170 742 14580 884
rect 9562 654 9986 712
rect 14170 704 14588 742
rect -14594 522 -14180 560
rect -11154 582 -11054 648
rect -9986 582 -9576 654
rect -14594 380 -14188 522
rect -11154 482 -9576 582
rect 9576 542 9986 654
rect 14180 560 14588 704
rect 9576 482 9994 542
rect 14180 522 14594 560
rect -14598 342 -14188 380
rect -9994 370 -9586 482
rect -14598 200 -14194 342
rect -9998 312 -9586 370
rect 9586 370 9994 482
rect 14188 380 14594 522
rect 9586 312 9998 370
rect 14188 342 14598 380
rect -9998 200 -9594 312
rect -14600 160 -14194 200
rect -14600 -160 -14198 160
rect -10000 142 -9594 200
rect 9594 200 9998 312
rect 14194 200 14598 342
rect 9594 142 10000 200
rect 14194 160 14600 200
rect -10000 -142 -9598 142
rect 9598 -142 10000 142
rect -14600 -198 -14194 -160
rect -10000 -198 -9594 -142
rect -14598 -342 -14194 -198
rect -9998 -312 -9594 -198
rect 9594 -200 10000 -142
rect 14198 -160 14600 160
rect 14194 -200 14600 -160
rect 9594 -312 9998 -200
rect -14598 -380 -14188 -342
rect -9998 -370 -9586 -312
rect -14594 -408 -14188 -380
rect -14594 -488 -12284 -408
rect -9994 -482 -9586 -370
rect 9586 -370 9998 -312
rect 14194 -342 14598 -200
rect 9586 -482 9994 -370
rect -14594 -522 -14188 -488
rect -14594 -560 -14180 -522
rect -9994 -542 -9576 -482
rect -14588 -704 -14180 -560
rect -9986 -654 -9576 -542
rect 9576 -542 9994 -482
rect 14188 -380 14598 -342
rect 14188 -522 14594 -380
rect 9576 -654 9986 -542
rect -14588 -742 -14170 -704
rect -9986 -712 -9562 -654
rect -14580 -884 -14170 -742
rect -9976 -824 -9562 -712
rect 9562 -712 9986 -654
rect 14180 -560 14594 -522
rect 14180 -704 14588 -560
rect 9562 -824 9976 -712
rect -9976 -882 -9546 -824
rect -14580 -922 -14158 -884
rect -14570 -1064 -14158 -922
rect -9962 -994 -9546 -882
rect 9546 -882 9976 -824
rect 14170 -742 14588 -704
rect 9546 -994 9962 -882
rect 14170 -884 14580 -742
rect -9962 -1054 -9526 -994
rect -14570 -1104 -14144 -1064
rect -14558 -1244 -14144 -1104
rect -9946 -1162 -9526 -1054
rect 9526 -1054 9962 -994
rect 14158 -922 14580 -884
rect 9526 -1140 9946 -1054
rect 14158 -1064 14570 -922
rect 14144 -1104 14570 -1064
rect 9526 -1162 11600 -1140
rect -9946 -1224 -9504 -1162
rect -14558 -1284 -14126 -1244
rect -14544 -1424 -14126 -1284
rect -9926 -1332 -9504 -1224
rect 9504 -1240 11600 -1162
rect 9504 -1332 9926 -1240
rect 14144 -1244 14558 -1104
rect -9926 -1394 -9478 -1332
rect -14544 -1464 -14108 -1424
rect -14526 -1604 -14108 -1464
rect -9904 -1500 -9478 -1394
rect 9478 -1394 9926 -1332
rect 14126 -1284 14558 -1244
rect 9478 -1500 9904 -1394
rect 14126 -1424 14544 -1284
rect -9904 -1562 -9450 -1500
rect -14526 -1644 -14086 -1604
rect -14508 -1784 -14086 -1644
rect -9878 -1668 -9450 -1562
rect 9450 -1562 9904 -1500
rect 14108 -1464 14544 -1424
rect 9450 -1668 9878 -1562
rect 14108 -1604 14526 -1464
rect -9878 -1732 -9418 -1668
rect -14508 -1824 -14062 -1784
rect -14486 -1962 -14062 -1824
rect -9850 -1836 -9418 -1732
rect 9418 -1732 9878 -1668
rect 14086 -1644 14526 -1604
rect 9418 -1836 9850 -1732
rect 14086 -1784 14508 -1644
rect -9850 -1900 -9384 -1836
rect -14486 -2004 -14036 -1962
rect -14462 -2140 -14036 -2004
rect -9818 -2004 -9384 -1900
rect 9384 -1900 9850 -1836
rect 14062 -1824 14508 -1784
rect 9384 -2004 9818 -1900
rect 14062 -1962 14486 -1824
rect -9818 -2068 -9348 -2004
rect -14462 -2184 -14008 -2140
rect -14436 -2320 -14008 -2184
rect -9784 -2170 -9348 -2068
rect 9348 -2068 9818 -2004
rect 14036 -2004 14486 -1962
rect 9348 -2170 9784 -2068
rect 14036 -2140 14462 -2004
rect 14008 -2156 14462 -2140
rect -9784 -2236 -9308 -2170
rect -14436 -2362 -13976 -2320
rect -14408 -2498 -13976 -2362
rect -9748 -2336 -9308 -2236
rect 9308 -2236 9784 -2170
rect 12196 -2184 14462 -2156
rect 12196 -2236 14436 -2184
rect 9308 -2336 9748 -2236
rect 14008 -2320 14436 -2236
rect -9748 -2404 -9266 -2336
rect -14408 -2540 -13944 -2498
rect -14376 -2674 -13944 -2540
rect -9708 -2500 -9266 -2404
rect 9266 -2404 9748 -2336
rect 13976 -2362 14436 -2320
rect 9266 -2500 9708 -2404
rect 13976 -2498 14408 -2362
rect -9708 -2570 -9220 -2500
rect -9666 -2664 -9220 -2570
rect 9220 -2570 9708 -2500
rect 13944 -2540 14408 -2498
rect 9220 -2664 9666 -2570
rect -14376 -2720 -13908 -2674
rect -14344 -2852 -13908 -2720
rect -9666 -2736 -9170 -2664
rect -9620 -2828 -9170 -2736
rect 9170 -2736 9666 -2664
rect 13944 -2674 14376 -2540
rect 13908 -2720 14376 -2674
rect 9170 -2828 9620 -2736
rect -14344 -2898 -13872 -2852
rect -14308 -3028 -13872 -2898
rect -9620 -2900 -9120 -2828
rect -14308 -3074 -13832 -3028
rect -14272 -3204 -13832 -3074
rect -12364 -3116 -12264 -2928
rect -9570 -2990 -9120 -2900
rect 9120 -2900 9620 -2828
rect 13908 -2852 14344 -2720
rect 13872 -2898 14344 -2852
rect 9120 -2990 9570 -2900
rect -9570 -3064 -9066 -2990
rect -9520 -3116 -9066 -3064
rect -12364 -3150 -9066 -3116
rect 9066 -3064 9570 -2990
rect 13872 -3028 14308 -2898
rect 9066 -3150 9520 -3064
rect -14272 -3252 -13790 -3204
rect -12364 -3216 -9008 -3150
rect -9520 -3228 -9008 -3216
rect -14232 -3380 -13790 -3252
rect -9466 -3312 -9008 -3228
rect 9008 -3228 9520 -3150
rect 13832 -3074 14308 -3028
rect 13832 -3204 14272 -3074
rect 9008 -3312 9466 -3228
rect -14232 -3428 -13746 -3380
rect -9466 -3390 -8948 -3312
rect -14190 -3556 -13746 -3428
rect -9408 -3470 -8948 -3390
rect 8948 -3390 9466 -3312
rect 13790 -3252 14272 -3204
rect 13790 -3380 14232 -3252
rect 8948 -3470 9408 -3390
rect -9408 -3550 -8886 -3470
rect -14190 -3604 -13700 -3556
rect -14146 -3660 -13700 -3604
rect -9348 -3628 -8886 -3550
rect 8886 -3550 9408 -3470
rect 13746 -3428 14232 -3380
rect 8886 -3628 9348 -3550
rect 13746 -3556 14190 -3428
rect -14146 -3740 -10000 -3660
rect -9348 -3712 -8820 -3628
rect -14146 -3780 -13652 -3740
rect -14100 -3904 -13652 -3780
rect -14100 -3956 -13602 -3904
rect -10080 -3906 -10000 -3740
rect -9286 -3786 -8820 -3712
rect 8820 -3712 9348 -3628
rect 13700 -3604 14190 -3556
rect 8820 -3786 9286 -3712
rect 13700 -3730 14146 -3604
rect -9286 -3870 -8752 -3786
rect -14052 -4076 -13602 -3956
rect -9220 -3940 -8752 -3870
rect 8752 -3870 9286 -3786
rect 13652 -3780 14146 -3730
rect 8752 -3940 9220 -3870
rect 13652 -3904 14100 -3780
rect -9220 -4028 -8680 -3940
rect -14052 -4130 -13550 -4076
rect -14002 -4248 -13550 -4130
rect -9152 -4096 -8680 -4028
rect 8680 -4028 9220 -3940
rect 13602 -3956 14100 -3904
rect 8680 -4096 9152 -4028
rect 13602 -4076 14052 -3956
rect -9152 -4186 -8608 -4096
rect -9080 -4248 -8608 -4186
rect 8608 -4186 9152 -4096
rect 13550 -4130 14052 -4076
rect 8608 -4248 9080 -4186
rect 13550 -4248 14002 -4130
rect -14002 -4304 -13494 -4248
rect -13950 -4420 -13494 -4304
rect -9080 -4340 -8530 -4248
rect -9008 -4400 -8530 -4340
rect 8530 -4340 9080 -4248
rect 13494 -4304 14002 -4248
rect 8530 -4400 9008 -4340
rect -13950 -4476 -13438 -4420
rect -13894 -4592 -13438 -4476
rect -9008 -4496 -8452 -4400
rect -8930 -4550 -8452 -4496
rect 8452 -4496 9008 -4400
rect 13494 -4420 13950 -4304
rect 13438 -4476 13950 -4420
rect 8452 -4550 8930 -4496
rect -13894 -4648 -13378 -4592
rect -8930 -4648 -8370 -4550
rect -13838 -4762 -13378 -4648
rect -8852 -4700 -8370 -4648
rect 8370 -4648 8930 -4550
rect 13438 -4592 13894 -4476
rect 13378 -4648 13894 -4592
rect 8370 -4700 8852 -4648
rect -13838 -4820 -13316 -4762
rect -8852 -4800 -8286 -4700
rect -13778 -4932 -13316 -4820
rect -8770 -4846 -8286 -4800
rect 8286 -4800 8852 -4700
rect 12176 -4776 12432 -4676
rect 13378 -4762 13838 -4648
rect 8286 -4846 8770 -4800
rect -13778 -4992 -13254 -4932
rect -8770 -4950 -8200 -4846
rect -13716 -5100 -13254 -4992
rect -8686 -4992 -8200 -4950
rect 8200 -4900 8770 -4846
rect 12332 -4900 12432 -4776
rect 8200 -4992 12432 -4900
rect 13316 -4820 13838 -4762
rect 13316 -4932 13778 -4820
rect -8686 -5100 -8110 -4992
rect -13716 -5162 -13188 -5100
rect -13654 -5268 -13188 -5162
rect -8600 -5136 -8110 -5100
rect 8110 -5000 12432 -4992
rect 13254 -4992 13778 -4932
rect 8110 -5100 8686 -5000
rect 13254 -5100 13716 -4992
rect 8110 -5136 8600 -5100
rect -8600 -5246 -8018 -5136
rect -13654 -5332 -13120 -5268
rect -13588 -5434 -13120 -5332
rect -8510 -5280 -8018 -5246
rect 8018 -5246 8600 -5136
rect 13188 -5162 13716 -5100
rect 8018 -5280 8510 -5246
rect 13188 -5268 13654 -5162
rect -8510 -5392 -7924 -5280
rect -8418 -5420 -7924 -5392
rect 7924 -5392 8510 -5280
rect 13120 -5332 13654 -5268
rect 13120 -5390 13588 -5332
rect 7924 -5420 8418 -5392
rect -13588 -5500 -13050 -5434
rect -13520 -5600 -13050 -5500
rect -8418 -5536 -7826 -5420
rect -8324 -5560 -7826 -5536
rect 7826 -5536 8418 -5420
rect 10644 -5470 13588 -5390
rect 13050 -5500 13588 -5470
rect 7826 -5560 8324 -5536
rect -13520 -5668 -12978 -5600
rect -13450 -5766 -12978 -5668
rect -8324 -5680 -7728 -5560
rect -8226 -5696 -7728 -5680
rect 7728 -5680 8324 -5560
rect 13050 -5600 13520 -5500
rect 12978 -5668 13520 -5600
rect 7728 -5696 8226 -5680
rect -13450 -5834 -12904 -5766
rect -8226 -5820 -7626 -5696
rect -13378 -5930 -12904 -5834
rect -8128 -5832 -7626 -5820
rect 7626 -5820 8226 -5696
rect 12978 -5766 13450 -5668
rect 7626 -5832 8128 -5820
rect -13378 -6000 -12828 -5930
rect -8128 -5960 -7522 -5832
rect -13304 -6094 -12828 -6000
rect -8026 -5966 -7522 -5960
rect 7522 -5960 8128 -5832
rect 12904 -5834 13450 -5766
rect 12904 -5930 13378 -5834
rect 7522 -5966 8026 -5960
rect -13304 -6166 -12750 -6094
rect -8026 -6096 -7416 -5966
rect -13228 -6256 -12750 -6166
rect -7922 -6098 -7416 -6096
rect 7416 -6096 8026 -5966
rect 12828 -6000 13378 -5930
rect 12828 -6094 13304 -6000
rect 7416 -6098 7922 -6096
rect -7922 -6228 -7306 -6098
rect 7306 -6228 7922 -6098
rect -7922 -6232 -7196 -6228
rect -13228 -6330 -12670 -6256
rect -13150 -6416 -12670 -6330
rect -7816 -6346 -7196 -6232
rect -10100 -6356 -7196 -6346
rect 7196 -6232 7922 -6228
rect 12750 -6166 13304 -6094
rect 7196 -6356 7816 -6232
rect 12750 -6256 13228 -6166
rect -13150 -6494 -12588 -6416
rect -10100 -6446 -7082 -6356
rect -13070 -6578 -12588 -6494
rect -13070 -6656 -12504 -6578
rect -12988 -6736 -12504 -6656
rect -12988 -6816 -12418 -6736
rect -12904 -6894 -12418 -6816
rect -12904 -6978 -12330 -6894
rect -8086 -6922 -7986 -6446
rect -7706 -6482 -7082 -6446
rect 7082 -6366 7816 -6356
rect 12670 -6330 13228 -6256
rect 7082 -6482 7706 -6366
rect 12670 -6416 13150 -6330
rect -7706 -6498 -6966 -6482
rect -7596 -6606 -6966 -6498
rect 6966 -6498 7706 -6482
rect 12588 -6494 13150 -6416
rect 6966 -6606 7596 -6498
rect 12588 -6578 13070 -6494
rect -7596 -6628 -6848 -6606
rect -7482 -6728 -6848 -6628
rect 6848 -6628 7596 -6606
rect 6848 -6728 7482 -6628
rect -7482 -6756 -6728 -6728
rect -7366 -6848 -6728 -6756
rect 6728 -6756 7482 -6728
rect 12504 -6656 13070 -6578
rect 12504 -6736 12988 -6656
rect 6728 -6806 7366 -6756
rect 6728 -6848 9352 -6806
rect -7366 -6882 -6606 -6848
rect -12818 -7052 -12330 -6978
rect -7248 -6966 -6606 -6882
rect 6606 -6906 9352 -6848
rect 12418 -6816 12988 -6736
rect 12418 -6894 12904 -6816
rect 6606 -6966 7248 -6906
rect -7248 -7006 -6482 -6966
rect -12818 -7136 -12240 -7052
rect -7128 -7082 -6482 -7006
rect 6482 -7006 7248 -6966
rect 6482 -7082 7128 -7006
rect -7128 -7128 -6356 -7082
rect -12730 -7206 -12240 -7136
rect -7006 -7196 -6356 -7128
rect 6356 -7128 7128 -7082
rect 6356 -7196 7006 -7128
rect -12730 -7294 -12148 -7206
rect -7006 -7248 -6228 -7196
rect -12640 -7362 -12148 -7294
rect -6962 -7306 -6228 -7248
rect 6228 -7248 7006 -7196
rect 6228 -7306 6882 -7248
rect -12640 -7452 -12054 -7362
rect -6962 -7366 -6098 -7306
rect -6962 -7370 -6862 -7366
rect -12548 -7514 -12054 -7452
rect -6756 -7416 -6098 -7366
rect 6098 -7366 6882 -7306
rect 6098 -7416 6756 -7366
rect -6756 -7482 -5966 -7416
rect -12548 -7606 -11958 -7514
rect -6628 -7522 -5966 -7482
rect 5966 -7482 6756 -7416
rect 5966 -7522 6628 -7482
rect -6628 -7596 -5832 -7522
rect -12454 -7668 -11958 -7606
rect -6498 -7626 -5832 -7596
rect 5832 -7596 6628 -7522
rect 5832 -7626 6498 -7596
rect -12454 -7762 -11860 -7668
rect -6498 -7706 -5696 -7626
rect -12358 -7818 -11860 -7762
rect -6366 -7728 -5696 -7706
rect 5696 -7706 6498 -7626
rect 5696 -7728 6366 -7706
rect -6366 -7816 -5560 -7728
rect -12358 -7914 -11760 -7818
rect -12260 -7968 -11760 -7914
rect -6232 -7826 -5560 -7816
rect 5560 -7816 6366 -7728
rect 5560 -7826 6232 -7816
rect -6232 -7922 -5420 -7826
rect -6096 -7924 -5420 -7922
rect 5420 -7922 6232 -7826
rect 5420 -7924 6096 -7922
rect -12260 -8068 -11658 -7968
rect -6096 -8018 -5280 -7924
rect 5280 -8018 6096 -7924
rect -6096 -8026 -5136 -8018
rect -12160 -8116 -11658 -8068
rect -5960 -8110 -5136 -8026
rect 5136 -8026 6096 -8018
rect 5136 -8110 5960 -8026
rect -12160 -8218 -11554 -8116
rect -5960 -8128 -4992 -8110
rect -12058 -8264 -11554 -8218
rect -5820 -8200 -4992 -8128
rect 4992 -8128 5960 -8110
rect 4992 -8200 5820 -8128
rect 8190 -8140 8290 -6906
rect 9252 -8072 9352 -6906
rect 12330 -6978 12904 -6894
rect 12330 -7052 12818 -6978
rect 12240 -7136 12818 -7052
rect 12240 -7206 12730 -7136
rect 12148 -7294 12730 -7206
rect 12148 -7362 12640 -7294
rect 12054 -7452 12640 -7362
rect 12054 -7514 12548 -7452
rect 11958 -7606 12548 -7514
rect 11958 -7668 12454 -7606
rect 11860 -7762 12454 -7668
rect 11860 -7818 12358 -7762
rect 10624 -8072 10724 -7898
rect 11760 -7914 12358 -7818
rect 11760 -7968 12260 -7914
rect 9252 -8172 10724 -8072
rect 11658 -8068 12260 -7968
rect 11658 -8116 12160 -8068
rect -5820 -8226 -4846 -8200
rect -12058 -8368 -11448 -8264
rect -5680 -8286 -4846 -8226
rect 4846 -8226 5820 -8200
rect 11554 -8218 12160 -8116
rect 4846 -8286 5680 -8226
rect 11554 -8264 12058 -8218
rect -5680 -8324 -4700 -8286
rect -11954 -8408 -11448 -8368
rect -5536 -8370 -4700 -8324
rect 4700 -8324 5680 -8286
rect 4700 -8370 5536 -8324
rect -11954 -8516 -11342 -8408
rect -5536 -8418 -4550 -8370
rect -5392 -8452 -4550 -8418
rect 4550 -8418 5536 -8370
rect 11448 -8368 12058 -8264
rect 11448 -8408 11954 -8368
rect 4550 -8452 5392 -8418
rect -5392 -8510 -4400 -8452
rect -11848 -8554 -11342 -8516
rect -5290 -8530 -4400 -8510
rect 4400 -8510 5392 -8452
rect 4400 -8530 5246 -8510
rect -11848 -8664 -11232 -8554
rect -11742 -8696 -11232 -8664
rect -5290 -8600 -4248 -8530
rect -11742 -8808 -11122 -8696
rect -11632 -8838 -11122 -8808
rect -11632 -8954 -11008 -8838
rect -11522 -8978 -11008 -8954
rect -11522 -9096 -10894 -8978
rect -11408 -9116 -10894 -9096
rect -11408 -9238 -10778 -9116
rect -5290 -9152 -5190 -8600
rect -5100 -8608 -4248 -8600
rect 4248 -8600 5246 -8530
rect 11342 -8516 11954 -8408
rect 11342 -8554 11848 -8516
rect 4248 -8608 5194 -8600
rect -5100 -8680 -4096 -8608
rect 4096 -8680 5194 -8608
rect -5100 -8686 -3940 -8680
rect -4950 -8752 -3940 -8686
rect 3940 -8686 5194 -8680
rect 3940 -8752 4950 -8686
rect -4950 -8770 -3786 -8752
rect -4800 -8820 -3786 -8770
rect 3786 -8770 4950 -8752
rect 3786 -8820 4800 -8770
rect -4800 -8852 -3628 -8820
rect -4648 -8886 -3628 -8852
rect 3628 -8852 4800 -8820
rect 3628 -8886 4648 -8852
rect -4648 -8930 -3470 -8886
rect -4496 -8948 -3470 -8930
rect 3470 -8930 4648 -8886
rect 3470 -8948 4496 -8930
rect -4496 -9008 -3312 -8948
rect 3312 -9008 4496 -8948
rect -4340 -9066 -3150 -9008
rect 3150 -9066 4340 -9008
rect -4340 -9080 -2990 -9066
rect -4186 -9120 -2990 -9080
rect 2990 -9080 4340 -9066
rect 2990 -9120 4186 -9080
rect -4186 -9152 -2828 -9120
rect -4028 -9170 -2828 -9152
rect 2828 -9152 4186 -9120
rect 2828 -9170 4028 -9152
rect -4028 -9220 -2664 -9170
rect 2664 -9220 4028 -9170
rect -11294 -9254 -10778 -9238
rect -11294 -9378 -10660 -9254
rect -3870 -9266 -2500 -9220
rect 2500 -9266 3870 -9220
rect -3870 -9286 -2336 -9266
rect -3712 -9308 -2336 -9286
rect 2336 -9286 3870 -9266
rect 2336 -9308 3712 -9286
rect -3712 -9348 -2170 -9308
rect 2170 -9348 3712 -9308
rect -11178 -9390 -10660 -9378
rect -11178 -9516 -10540 -9390
rect -11060 -9524 -10540 -9516
rect -11060 -9654 -10420 -9524
rect -10940 -9656 -10420 -9654
rect -10940 -9788 -10296 -9656
rect -10940 -9790 -10172 -9788
rect -10820 -9918 -10172 -9790
rect -10820 -9924 -10046 -9918
rect -10696 -10046 -10046 -9924
rect -10696 -10056 -9918 -10046
rect -10572 -10172 -9918 -10056
rect -10572 -10188 -9788 -10172
rect -10446 -10296 -9788 -10188
rect -10446 -10318 -9656 -10296
rect -10318 -10420 -9656 -10318
rect -10318 -10446 -9524 -10420
rect -10188 -10540 -9524 -10446
rect -10188 -10572 -9390 -10540
rect -10056 -10660 -9390 -10572
rect -10056 -10696 -9254 -10660
rect -9924 -10778 -9254 -10696
rect -9924 -10820 -9116 -10778
rect -9790 -10894 -9116 -10820
rect -9790 -10940 -8978 -10894
rect -9654 -11008 -8978 -10940
rect -9654 -11060 -8838 -11008
rect -9516 -11122 -8838 -11060
rect -9516 -11178 -8696 -11122
rect -9378 -11232 -8696 -11178
rect -9378 -11294 -8554 -11232
rect -9238 -11342 -8554 -11294
rect -9238 -11408 -8408 -11342
rect -9096 -11448 -8408 -11408
rect -9096 -11522 -8264 -11448
rect -8954 -11554 -8264 -11522
rect -8954 -11632 -8116 -11554
rect -8808 -11658 -8116 -11632
rect -8066 -11658 -7986 -9362
rect -3550 -9384 -2004 -9348
rect 2004 -9384 3550 -9348
rect -3550 -9408 -1836 -9384
rect -3390 -9418 -1836 -9408
rect 1836 -9408 3550 -9384
rect 1836 -9418 3390 -9408
rect -3390 -9450 -1668 -9418
rect 1668 -9450 3390 -9418
rect -3390 -9466 -1500 -9450
rect -3228 -9478 -1500 -9466
rect 1500 -9466 3390 -9450
rect 1500 -9478 3228 -9466
rect -3228 -9504 -1332 -9478
rect 1332 -9504 3228 -9478
rect -3228 -9520 -1162 -9504
rect -3064 -9526 -1162 -9520
rect 1162 -9520 3228 -9504
rect 1162 -9526 3064 -9520
rect -3064 -9546 -994 -9526
rect 994 -9546 3064 -9526
rect -3064 -9562 -824 -9546
rect 824 -9562 3064 -9546
rect -3064 -9570 -654 -9562
rect -2900 -9576 -654 -9570
rect 654 -9570 3064 -9562
rect 654 -9576 2900 -9570
rect -2900 -9586 -482 -9576
rect 482 -9586 2900 -9576
rect -2900 -9594 -312 -9586
rect 312 -9594 2900 -9586
rect -2900 -9598 -142 -9594
rect 142 -9598 2900 -9594
rect -2900 -9620 2900 -9598
rect -2736 -9666 2736 -9620
rect -2570 -9708 2570 -9666
rect -2404 -9748 2404 -9708
rect -2236 -9784 2236 -9748
rect -2068 -9818 2068 -9784
rect -1960 -9850 1900 -9818
rect -1960 -10458 -1860 -9850
rect -1732 -9878 1732 -9850
rect -1562 -9904 1562 -9878
rect -1394 -9926 1394 -9904
rect -1224 -9946 1224 -9926
rect -1054 -9962 1054 -9946
rect -882 -9976 882 -9962
rect -712 -9986 712 -9976
rect -542 -9994 542 -9986
rect -370 -9998 370 -9994
rect -200 -10000 198 -9998
rect 1606 -10726 1706 -9878
rect 5094 -9930 5194 -8686
rect 11232 -8664 11848 -8554
rect 11232 -8696 11742 -8664
rect 11122 -8808 11742 -8696
rect 11122 -8838 11632 -8808
rect 11008 -8954 11632 -8838
rect 11008 -8978 11522 -8954
rect 10894 -9096 11522 -8978
rect 10894 -9116 11408 -9096
rect 10778 -9238 11408 -9116
rect 10778 -9254 11294 -9238
rect 10660 -9378 11294 -9254
rect 10660 -9390 11178 -9378
rect 10540 -9516 11178 -9390
rect 10540 -9524 11060 -9516
rect 10420 -9654 11060 -9524
rect 10420 -9656 10940 -9654
rect 10296 -9788 10940 -9656
rect 10172 -9790 10940 -9788
rect 10172 -9918 10820 -9790
rect 10046 -9924 10820 -9918
rect 10046 -10046 10696 -9924
rect 9918 -10056 10696 -10046
rect 9918 -10172 10572 -10056
rect 9788 -10188 10572 -10172
rect 9788 -10296 10446 -10188
rect 9656 -10318 10446 -10296
rect 9656 -10420 10318 -10318
rect 9524 -10446 10318 -10420
rect 9524 -10540 10188 -10446
rect 9390 -10572 10188 -10540
rect 8210 -11448 8290 -10580
rect 9390 -10660 10056 -10572
rect 9254 -10696 10056 -10660
rect 9254 -10778 9924 -10696
rect 9116 -10820 9924 -10778
rect 9116 -10894 9790 -10820
rect 8978 -10940 9790 -10894
rect 8978 -11008 9654 -10940
rect 8838 -11060 9654 -11008
rect 8838 -11122 9516 -11060
rect 8696 -11178 9516 -11122
rect 8696 -11232 9378 -11178
rect 8554 -11294 9378 -11232
rect 8554 -11342 9238 -11294
rect 8408 -11408 9238 -11342
rect 8408 -11448 9096 -11408
rect 8210 -11522 9096 -11448
rect 8210 -11554 8954 -11522
rect -8808 -11742 -7968 -11658
rect -8664 -11760 -7968 -11742
rect -8664 -11848 -7818 -11760
rect -8516 -11860 -7818 -11848
rect -8516 -11954 -7668 -11860
rect -8368 -11958 -7668 -11954
rect -8368 -12054 -7514 -11958
rect -8368 -12058 -7362 -12054
rect -8218 -12148 -7362 -12058
rect -8218 -12160 -7206 -12148
rect -8068 -12240 -7206 -12160
rect -8068 -12260 -7052 -12240
rect -7914 -12330 -7052 -12260
rect -7914 -12358 -6894 -12330
rect -7762 -12418 -6894 -12358
rect -7762 -12454 -6736 -12418
rect -7606 -12504 -6736 -12454
rect -7606 -12548 -6578 -12504
rect -7452 -12588 -6578 -12548
rect -7452 -12640 -6416 -12588
rect -7294 -12670 -6416 -12640
rect -7294 -12730 -6256 -12670
rect -7136 -12750 -6256 -12730
rect -7136 -12818 -6094 -12750
rect -6978 -12828 -6094 -12818
rect -6978 -12904 -5930 -12828
rect -6816 -12978 -5766 -12904
rect -6816 -12988 -5600 -12978
rect -6656 -13050 -5600 -12988
rect -6656 -13070 -5434 -13050
rect -6494 -13120 -5434 -13070
rect -5270 -13120 -5190 -11592
rect 8116 -11632 8954 -11554
rect 8116 -11658 8808 -11632
rect 7968 -11742 8808 -11658
rect 7968 -11760 8664 -11742
rect 7818 -11848 8664 -11760
rect 7818 -11860 8516 -11848
rect 7668 -11954 8516 -11860
rect 7668 -11958 8368 -11954
rect 7514 -12054 8368 -11958
rect 7362 -12058 8368 -12054
rect 7362 -12148 8218 -12058
rect 7206 -12160 8218 -12148
rect 7206 -12240 8068 -12160
rect 7052 -12260 8068 -12240
rect 7052 -12330 7914 -12260
rect 6894 -12358 7914 -12330
rect -6494 -13150 -5190 -13120
rect -6330 -13188 -5190 -13150
rect -6330 -13228 -5100 -13188
rect -6166 -13254 -5100 -13228
rect -6166 -13304 -4932 -13254
rect -6000 -13316 -4932 -13304
rect -6000 -13378 -4762 -13316
rect -1940 -13368 -1860 -12898
rect -5834 -13438 -4592 -13378
rect -5834 -13450 -4420 -13438
rect -5668 -13494 -4420 -13450
rect -1982 -13448 -1860 -13368
rect -5668 -13520 -4248 -13494
rect -5500 -13550 -4248 -13520
rect -5500 -13588 -4076 -13550
rect -5332 -13602 -4076 -13588
rect -5332 -13652 -3904 -13602
rect -5332 -13654 -3730 -13652
rect -5162 -13700 -3730 -13654
rect -5162 -13716 -3556 -13700
rect -4992 -13746 -3556 -13716
rect -4992 -13778 -3380 -13746
rect -4820 -13790 -3380 -13778
rect -4820 -13832 -3204 -13790
rect -4820 -13838 -3028 -13832
rect -4648 -13872 -3028 -13838
rect -4648 -13894 -2852 -13872
rect -4476 -13908 -2852 -13894
rect -4476 -13944 -2674 -13908
rect -4476 -13950 -2498 -13944
rect -4304 -13976 -2498 -13950
rect -4304 -14002 -2320 -13976
rect -4130 -14008 -2320 -14002
rect -4130 -14036 -2140 -14008
rect -1982 -14036 -1902 -13448
rect -4130 -14052 -1902 -14036
rect -3956 -14062 -1902 -14052
rect -3956 -14086 -1784 -14062
rect 1626 -14086 1706 -13166
rect 5114 -13188 5194 -12370
rect 6894 -12418 7762 -12358
rect 6736 -12454 7762 -12418
rect 6736 -12504 7606 -12454
rect 6578 -12548 7606 -12504
rect 6578 -12588 7452 -12548
rect 6416 -12640 7452 -12588
rect 6416 -12670 7294 -12640
rect 6256 -12730 7294 -12670
rect 6256 -12750 7136 -12730
rect 6094 -12818 7136 -12750
rect 6094 -12828 6978 -12818
rect 5930 -12904 6978 -12828
rect 5766 -12978 6816 -12904
rect 5600 -12988 6816 -12978
rect 5600 -13050 6656 -12988
rect 5434 -13070 6656 -13050
rect 5434 -13120 6494 -13070
rect 5268 -13150 6494 -13120
rect 5268 -13188 6330 -13150
rect 5100 -13228 6330 -13188
rect 5100 -13254 6166 -13228
rect 4932 -13304 6166 -13254
rect 4932 -13316 6000 -13304
rect 4762 -13378 6000 -13316
rect 4592 -13438 5834 -13378
rect 4420 -13450 5834 -13438
rect 4420 -13494 5668 -13450
rect 4248 -13520 5668 -13494
rect 4248 -13550 5500 -13520
rect 4076 -13588 5500 -13550
rect 4076 -13602 5332 -13588
rect 3904 -13652 5332 -13602
rect 3730 -13654 5332 -13652
rect 3730 -13700 5162 -13654
rect 3556 -13716 5162 -13700
rect 3556 -13746 4992 -13716
rect 3380 -13778 4992 -13746
rect 3380 -13790 4820 -13778
rect 3204 -13832 4820 -13790
rect 3028 -13838 4820 -13832
rect 3028 -13872 4648 -13838
rect 2852 -13894 4648 -13872
rect 2852 -13908 4476 -13894
rect 2674 -13944 4476 -13908
rect 2498 -13950 4476 -13944
rect 2498 -13976 4304 -13950
rect 2320 -14002 4304 -13976
rect 2320 -14008 4130 -14002
rect 2140 -14036 4130 -14008
rect 1962 -14052 4130 -14036
rect 1962 -14062 3956 -14052
rect 1784 -14086 3956 -14062
rect -3956 -14100 -1604 -14086
rect -3780 -14108 -1604 -14100
rect 1604 -14100 3956 -14086
rect 1604 -14108 3780 -14100
rect -3780 -14126 -1424 -14108
rect 1424 -14126 3780 -14108
rect -3780 -14144 -1244 -14126
rect 1244 -14144 3780 -14126
rect -3780 -14146 -1064 -14144
rect -3604 -14158 -1064 -14146
rect 1064 -14146 3780 -14144
rect 1064 -14158 3604 -14146
rect -3604 -14170 -884 -14158
rect 884 -14170 3604 -14158
rect -3604 -14180 -704 -14170
rect 704 -14180 3604 -14170
rect -3604 -14188 -522 -14180
rect 522 -14188 3604 -14180
rect -3604 -14190 -342 -14188
rect -3428 -14194 -342 -14190
rect 342 -14190 3604 -14188
rect 342 -14194 3428 -14190
rect -3428 -14198 -160 -14194
rect 160 -14198 3428 -14194
rect -3428 -14232 3428 -14198
rect -3252 -14272 3252 -14232
rect -3074 -14308 3074 -14272
rect -2898 -14344 2898 -14308
rect -2720 -14376 2720 -14344
rect -2540 -14408 2540 -14376
rect -2362 -14436 2362 -14408
rect -2184 -14462 2184 -14436
rect -2004 -14486 2004 -14462
rect -1824 -14508 1824 -14486
rect -1644 -14526 1644 -14508
rect -1464 -14544 1464 -14526
rect -1284 -14558 1284 -14544
rect -1104 -14570 1104 -14558
rect -922 -14580 922 -14570
rect -742 -14588 742 -14580
rect -560 -14594 560 -14588
rect -380 -14598 380 -14594
rect -200 -14600 198 -14598
use skullfet_inverter  skullfet_inverter_0
timestamp 1712756528
transform 1 0 11000 0 1 -1400
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_1
timestamp 1712756528
transform -1 0 12776 0 1 2136
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_2
timestamp 1712756528
transform 1 0 8914 0 1 5358
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_3
timestamp 1712756528
transform 1 0 6480 0 1 7980
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_4
timestamp 1712756528
transform 1 0 3384 0 1 9770
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_5
timestamp 1712756528
transform 1 0 -104 0 1 10566
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_6
timestamp 1712756528
transform 1 0 -3670 0 1 10298
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_7
timestamp 1712756528
transform 1 0 -6998 0 1 8992
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_8
timestamp 1712756528
transform 1 0 -9796 0 1 6762
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_9
timestamp 1712756528
transform 1 0 -11810 0 1 3806
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_10
timestamp 1712756528
transform -1 0 -10554 0 1 388
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_11
timestamp 1712756528
transform 1 0 -12864 0 1 -3188
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_12
timestamp 1712756528
transform -1 0 -9500 0 1 -6606
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_13
timestamp 1712756528
transform -1 0 -7486 0 -1 -6662
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_14
timestamp 1712756528
transform -1 0 -4690 0 -1 -8892
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_15
timestamp 1712756528
transform -1 0 -1360 0 -1 -10198
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_16
timestamp 1712756528
transform -1 0 2206 0 -1 -10466
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_17
timestamp 1712756528
transform -1 0 5694 0 -1 -9670
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_18
timestamp 1712756528
transform -1 0 8790 0 -1 -7880
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_19
timestamp 1712756528
transform -1 0 11224 0 1 -8158
box 410 120 1900 2780
use skullfet_inverter  skullfet_inverter_20
timestamp 1712756528
transform -1 0 12776 0 1 -4936
box 410 120 1900 2780
<< end >>
