* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5]
+ uo_out[6] uo_out[7] uo_out[0] VPWR VGND
X0 VGND.t35 uo_out[0].t2 ring_0/skullfet_inverter_6.A VGND.t34 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X1 VGND.t39 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t38 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X2 ring_0/skullfet_inverter_6.A uo_out[0].t3 VPWR.t35 VPWR.t34 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X3 VGND.t11 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VGND.t10 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X4 VGND.t5 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t4 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X5 VGND.t25 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_8.A VGND.t24 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X6 VGND.t23 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t22 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X7 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VPWR.t39 VPWR.t38 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X8 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t29 VGND.t28 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X9 VGND.t33 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t32 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X10 VGND.t17 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t16 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X11 VPWR.t15 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VPWR.t14 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X12 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t31 VGND.t30 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X13 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_7.A VPWR.t25 VPWR.t24 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X14 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_8.A VPWR.t3 VPWR.t2 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X15 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VPWR.t33 VPWR.t32 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X16 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VPWR.t23 VPWR.t22 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X17 VGND.t21 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t20 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X18 VPWR.t37 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VPWR.t36 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X19 VPWR.t19 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VPWR.t18 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X20 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VPWR.t17 VPWR.t16 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X21 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X22 VPWR.t29 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VPWR.t28 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X23 VGND.t7 ring_0/skullfet_inverter_4.A uo_out[0].t0 VGND.t6 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X24 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VPWR.t13 VPWR.t12 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X25 VGND.t41 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t40 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X26 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VPWR.t21 VPWR.t20 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X27 VPWR.t1 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VPWR.t0 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X28 VGND.t9 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t8 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X29 uo_out[0].t1 ring_0/skullfet_inverter_4.A VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X30 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VPWR.t41 VPWR.t40 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X31 VGND.t13 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t12 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X32 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VPWR.t9 VPWR.t8 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X33 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VPWR.t27 VPWR.t26 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X34 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X35 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X36 VPWR.t31 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VPWR.t30 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X37 VGND.t27 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VGND.t26 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X38 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t37 VGND.t36 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X39 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t19 VGND.t18 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X40 VGND.t3 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_9.A VGND.t2 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X41 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VPWR.t5 VPWR.t4 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
R0 uo_out[0] uo_out[0].t1 984.356
R1 uo_out[0].n0 uo_out[0].t2 582.378
R2 uo_out[0].n1 uo_out[0].t3 566.953
R3 uo_out[0].n4 uo_out[0].t0 478.87
R4 uo_out[0].n1 uo_out[0].n0 424.161
R5 uo_out[0].n2 uo_out[0].n0 204.481
R6 uo_out[0] uo_out[0].n1 201.921
R7 uo_out[0].n3 uo_out[0] 19.3513
R8 uo_out[0].n2 uo_out[0] 10.2405
R9 uo_out[0] uo_out[0].n4 10.2405
R10 uo_out[0].n4 uo_out[0].n3 7.5409
R11 uo_out[0].n3 uo_out[0].n2 5.01603
R12 VGND.n305 VGND.n62 171881
R13 VGND.n323 VGND.n322 156689
R14 VGND.n65 VGND.t22 151322
R15 VGND.n302 VGND.n97 130569
R16 VGND.n349 VGND.n348 130542
R17 VGND.n149 VGND.n3 48636.9
R18 VGND.n308 VGND.n97 45450.3
R19 VGND.n350 VGND.n349 44132.5
R20 VGND.n302 VGND.n301 44106
R21 VGND.n303 VGND.n99 43377.2
R22 VGND.n301 VGND.n300 30151.8
R23 VGND.n351 VGND.n350 30151.8
R24 VGND.n301 VGND.n100 29891.4
R25 VGND.n350 VGND.n1 29891.4
R26 VGND.n308 VGND.n62 16600.2
R27 VGND.n159 VGND.n154 16072.7
R28 VGND.n98 VGND.n61 14081.5
R29 VGND.n144 VGND.n143 12272.6
R30 VGND.n167 VGND.n144 12077.4
R31 VGND.n309 VGND.n308 11373.6
R32 VGND.n303 VGND.n302 10649.3
R33 VGND.n349 VGND.n3 10649.2
R34 VGND.n146 VGND.n144 6135.59
R35 VGND.n304 VGND.n303 6127.89
R36 VGND.t16 VGND.n158 4169.04
R37 VGND.n308 VGND.n96 3998.58
R38 VGND.n322 VGND.n321 3462.51
R39 VGND.n158 VGND.n157 3164.24
R40 VGND.n160 VGND.n159 3164.24
R41 VGND.n159 VGND.n156 3154.4
R42 VGND.n146 VGND.n145 3108.35
R43 VGND.n149 VGND.n146 3022.83
R44 VGND.n158 VGND.n154 2949.38
R45 VGND.n143 VGND.n98 2758.39
R46 VGND.n308 VGND.n307 2554.5
R47 VGND.n321 VGND.t40 2387.95
R48 VGND.n168 VGND.n98 2252.33
R49 VGND.n308 VGND.n304 2096.68
R50 VGND.n323 VGND.n62 1821.62
R51 VGND.n148 VGND.t36 1524.56
R52 VGND.n175 VGND.n99 1397.72
R53 VGND.n150 VGND.n149 1261.32
R54 VGND.n299 VGND.n298 1170
R55 VGND.n218 VGND.n95 1170
R56 VGND.n239 VGND.n96 1170
R57 VGND.n315 VGND.n64 1170
R58 VGND.n89 VGND.n63 1170
R59 VGND.n320 VGND.n319 1170
R60 VGND.n307 VGND.n306 1170
R61 VGND.n325 VGND.n324 1170
R62 VGND.n311 VGND.n310 1170
R63 VGND.n121 VGND.n120 1170
R64 VGND.n171 VGND.n170 1170
R65 VGND.n166 VGND.n165 1170
R66 VGND.n156 VGND.n155 1170
R67 VGND.n148 VGND.n147 1170
R68 VGND.n347 VGND.n346 1170
R69 VGND.n24 VGND.n2 1170
R70 VGND.n151 VGND.n150 1170
R71 VGND.n353 VGND.n352 1170
R72 VGND.n347 VGND.t28 1134.17
R73 VGND.t6 VGND.n99 1084.29
R74 VGND.n169 VGND.n168 1052.01
R75 VGND.n142 VGND.t8 1007.36
R76 VGND.t0 VGND.n323 876.702
R77 VGND.n97 VGND.t24 844.357
R78 VGND.n61 VGND.n4 843.24
R79 VGND.t18 VGND.n351 753.322
R80 VGND.n300 VGND.t20 733.058
R81 VGND.t22 VGND.n63 713.466
R82 VGND.t34 VGND.n100 698.659
R83 VGND.t14 VGND.n1 696.106
R84 VGND.n169 VGND.n142 637.375
R85 VGND.n321 VGND.n64 634.212
R86 VGND.n351 VGND.n2 585.742
R87 VGND.n300 VGND.n299 575.707
R88 VGND.n308 VGND.n95 546.717
R89 VGND.n352 VGND.n1 546.058
R90 VGND.n120 VGND.n100 531.929
R91 VGND.t40 VGND.n320 508.485
R92 VGND.n310 VGND.n309 333.548
R93 VGND.n154 VGND.t4 302.156
R94 VGND.n353 VGND.t19 282.339
R95 VGND.n24 VGND.t29 282.339
R96 VGND.n346 VGND.t31 282.339
R97 VGND.n325 VGND.t1 282.339
R98 VGND.n306 VGND.t39 282.339
R99 VGND.n155 VGND.t33 282.339
R100 VGND.n165 VGND.t11 282.339
R101 VGND.n147 VGND.t37 282.339
R102 VGND.n151 VGND.t15 282.339
R103 VGND.n157 VGND.t27 282.339
R104 VGND.n319 VGND.t41 282.339
R105 VGND.n218 VGND.t21 282.339
R106 VGND.n121 VGND.t7 282.339
R107 VGND.n171 VGND.t5 282.339
R108 VGND.n160 VGND.t17 282.339
R109 VGND.n175 VGND.t9 282.339
R110 VGND.n298 VGND.t35 282.339
R111 VGND.n239 VGND.t25 282.339
R112 VGND.n311 VGND.t3 282.339
R113 VGND.n315 VGND.t13 282.339
R114 VGND.n89 VGND.t23 282.339
R115 VGND.t24 VGND.n96 266.457
R116 VGND.t38 VGND.n305 248.936
R117 VGND.n158 VGND.t26 236.923
R118 VGND.n149 VGND.n148 212.281
R119 VGND.n166 VGND.n145 204.773
R120 VGND.n320 VGND.n65 190.542
R121 VGND.n307 VGND.t38 187.446
R122 VGND.n167 VGND.t10 183.096
R123 VGND.n352 VGND.t18 170.459
R124 VGND.n299 VGND.t34 167.052
R125 VGND.t28 VGND.n2 166.094
R126 VGND.t20 VGND.n95 162.857
R127 VGND.n308 VGND.t2 159.488
R128 VGND.n150 VGND.t14 158.115
R129 VGND.n120 VGND.t6 155.179
R130 VGND.n322 VGND.n63 144.5
R131 VGND.t10 VGND.n166 140.434
R132 VGND.n309 VGND.t12 132.02
R133 VGND.n324 VGND.t0 124.144
R134 VGND.n310 VGND.t2 122.326
R135 VGND.t32 VGND.n154 120.314
R136 VGND.n142 VGND.n99 112.184
R137 VGND.n170 VGND.t4 111.326
R138 VGND.n168 VGND.n167 104.849
R139 VGND.t12 VGND.n64 101.258
R140 VGND.n348 VGND.n4 100.996
R141 VGND.n156 VGND.t32 92.2804
R142 VGND.n159 VGND.t16 55.9751
R143 VGND.n348 VGND.n347 46.6396
R144 VGND.n143 VGND.n3 45.2738
R145 VGND.n324 VGND.n61 40.8576
R146 VGND.n170 VGND.n169 36.639
R147 VGND.n164 VGND.n153 20.9265
R148 VGND.n154 VGND.n145 20.0607
R149 VGND.n327 VGND.n60 17.0502
R150 VGND.n304 VGND.n98 14.7835
R151 VGND.n219 VGND.n218 13.3141
R152 VGND.n122 VGND.n121 13.3141
R153 VGND.n172 VGND.n171 13.3141
R154 VGND.n161 VGND.n160 13.3141
R155 VGND.n176 VGND.n175 13.3141
R156 VGND.n298 VGND.n297 13.3141
R157 VGND.n240 VGND.n239 13.3141
R158 VGND.n312 VGND.n311 13.3141
R159 VGND.n316 VGND.n315 13.3141
R160 VGND.n90 VGND.n89 13.3141
R161 VGND VGND.n24 13.2586
R162 VGND.n346 VGND 13.2586
R163 VGND VGND.n325 13.2586
R164 VGND.n306 VGND 13.2586
R165 VGND.n155 VGND 13.2586
R166 VGND.n165 VGND 13.2586
R167 VGND.n147 VGND 13.2586
R168 VGND VGND.n151 13.2586
R169 VGND.n157 VGND 13.2586
R170 VGND.n319 VGND 13.2586
R171 VGND VGND.n353 13.2586
R172 VGND VGND.n60 10.8878
R173 VGND.n317 VGND.n314 9.52816
R174 VGND VGND.n318 9.46719
R175 VGND.n162 VGND.n161 9.16992
R176 VGND VGND.n164 8.69654
R177 VGND.n173 VGND.n172 8.60727
R178 VGND.n326 VGND 8.50779
R179 VGND.n174 VGND.n173 8.47796
R180 VGND.n91 VGND.n90 7.73586
R181 VGND.n163 VGND 7.66873
R182 VGND VGND.n345 7.24133
R183 VGND.n177 VGND.n176 7.18609
R184 VGND.n317 VGND.n316 6.8256
R185 VGND VGND.n141 6.67637
R186 VGND.n313 VGND.n312 6.61112
R187 VGND.n196 VGND.n122 6.60276
R188 VGND.n25 VGND 6.5915
R189 VGND VGND.n0 6.55995
R190 VGND.n153 VGND 6.30778
R191 VGND.n273 VGND.n240 6.21471
R192 VGND.n152 VGND 6.20286
R193 VGND.n297 VGND.n296 6.13644
R194 VGND.n220 VGND.n219 5.99894
R195 VGND.n88 VGND.n87 3.93283
R196 VGND.n173 VGND.n141 3.52873
R197 VGND.n88 VGND 3.40017
R198 VGND.n153 VGND.n152 2.92676
R199 VGND.n318 VGND.n317 2.38171
R200 VGND.n305 VGND.n65 2.10058
R201 VGND.n4 VGND.t30 1.91332
R202 VGND.n164 VGND.n163 1.59945
R203 VGND.n152 VGND.n0 1.28972
R204 VGND.n92 VGND.n88 1.1273
R205 VGND.n163 VGND.n162 1.05629
R206 VGND.n318 VGND.n92 0.953601
R207 VGND.n162 VGND.n141 0.951859
R208 VGND.n66 uo_out[1] 0.8465
R209 VGND.n91 VGND.n60 0.753637
R210 VGND.n26 VGND.n0 0.663554
R211 VGND.n72 VGND.n71 0.5786
R212 VGND.n67 VGND.n66 0.577033
R213 VGND.n68 VGND.n67 0.577033
R214 VGND.n69 VGND.n68 0.577033
R215 VGND.n70 VGND.n69 0.577033
R216 VGND.n71 VGND.n70 0.577033
R217 VGND.n74 VGND.n73 0.577033
R218 VGND.n75 VGND.n74 0.577033
R219 VGND.n76 VGND.n75 0.577033
R220 VGND.n77 VGND.n76 0.577033
R221 VGND.n78 VGND.n77 0.577033
R222 VGND.n79 VGND.n78 0.577033
R223 VGND.n80 VGND.n79 0.577033
R224 VGND.n81 VGND.n80 0.577033
R225 VGND.n82 VGND.n81 0.577033
R226 VGND.n83 VGND.n82 0.577033
R227 VGND.n84 VGND.n83 0.577033
R228 VGND.n85 VGND.n84 0.577033
R229 VGND.n86 VGND.n85 0.577033
R230 VGND.n87 VGND.n86 0.577033
R231 VGND.n73 VGND.n72 0.575467
R232 VGND.n295 VGND.n294 0.457033
R233 VGND.n296 VGND.n101 0.297375
R234 VGND.n87 uio_oe[7] 0.2684
R235 VGND.n66 uo_out[2] 0.2684
R236 VGND.n67 uo_out[3] 0.2684
R237 VGND.n68 uo_out[4] 0.2684
R238 VGND.n69 uo_out[5] 0.2684
R239 VGND.n70 uo_out[6] 0.2684
R240 VGND.n71 uo_out[7] 0.2684
R241 VGND.n72 uio_out[0] 0.2684
R242 VGND.n73 uio_out[1] 0.2684
R243 VGND.n74 uio_out[2] 0.2684
R244 VGND.n75 uio_out[3] 0.2684
R245 VGND.n76 uio_out[4] 0.2684
R246 VGND.n77 uio_out[5] 0.2684
R247 VGND.n78 uio_out[6] 0.2684
R248 VGND.n79 uio_out[7] 0.2684
R249 VGND.n80 uio_oe[0] 0.2684
R250 VGND.n81 uio_oe[1] 0.2684
R251 VGND.n82 uio_oe[2] 0.2684
R252 VGND.n83 uio_oe[3] 0.2684
R253 VGND.n84 uio_oe[4] 0.2684
R254 VGND.n85 uio_oe[5] 0.2684
R255 VGND.n86 uio_oe[6] 0.2684
R256 VGND.n215 VGND.n101 0.240747
R257 VGND.n43 VGND.n7 0.232444
R258 VGND.n215 VGND.n214 0.201889
R259 VGND.n214 VGND.n213 0.183192
R260 VGND.n314 VGND.n93 0.181207
R261 VGND.n27 VGND.n26 0.177735
R262 VGND.n177 VGND.n174 0.15732
R263 VGND.n328 VGND.n327 0.155253
R264 VGND.n44 VGND.n43 0.152388
R265 VGND.n212 VGND.n211 0.145639
R266 VGND.n273 VGND.n272 0.14536
R267 VGND.n213 VGND.n212 0.14425
R268 VGND.n216 VGND.n215 0.135917
R269 VGND.n217 VGND.n101 0.135115
R270 VGND.n213 VGND.n103 0.134528
R271 VGND.n214 VGND.n102 0.133742
R272 VGND.n296 VGND.n295 0.133539
R273 VGND.n211 VGND.n105 0.133139
R274 VGND.n212 VGND.n104 0.133139
R275 VGND.n210 VGND.n106 0.13175
R276 VGND.n28 VGND.n22 0.131182
R277 VGND.n207 VGND.n109 0.131118
R278 VGND.n209 VGND.n107 0.131056
R279 VGND.n208 VGND.n108 0.130361
R280 VGND.n203 VGND.n113 0.129761
R281 VGND.n30 VGND.n20 0.129761
R282 VGND.n206 VGND.n110 0.129713
R283 VGND.n27 VGND.n23 0.129713
R284 VGND.n31 VGND.n19 0.128341
R285 VGND.n204 VGND.n112 0.128309
R286 VGND.n29 VGND.n21 0.128309
R287 VGND.n205 VGND.n111 0.128278
R288 VGND.n36 VGND.n14 0.12768
R289 VGND.n34 VGND.n16 0.127655
R290 VGND.n293 VGND.n292 0.127631
R291 VGND.n201 VGND.n115 0.127631
R292 VGND.n32 VGND.n18 0.127631
R293 VGND.n37 VGND.n13 0.126953
R294 VGND.n35 VGND.n15 0.126937
R295 VGND.n291 VGND.n221 0.12692
R296 VGND.n200 VGND.n116 0.12692
R297 VGND.n33 VGND.n17 0.12692
R298 VGND.n202 VGND.n114 0.126904
R299 VGND.n259 VGND.n254 0.126368
R300 VGND.n328 VGND.n59 0.126345
R301 VGND.n330 VGND.n57 0.126333
R302 VGND.n332 VGND.n55 0.126322
R303 VGND.n334 VGND.n53 0.126312
R304 VGND.n42 VGND.n8 0.126244
R305 VGND.n288 VGND.n224 0.126218
R306 VGND.n197 VGND.n119 0.126218
R307 VGND.n290 VGND.n222 0.12621
R308 VGND.n199 VGND.n117 0.12621
R309 VGND.n285 VGND.n227 0.1255
R310 VGND.n286 VGND.n226 0.1255
R311 VGND.n287 VGND.n225 0.1255
R312 VGND.n289 VGND.n223 0.1255
R313 VGND.n193 VGND.n125 0.1255
R314 VGND.n194 VGND.n124 0.1255
R315 VGND.n195 VGND.n123 0.1255
R316 VGND.n198 VGND.n118 0.1255
R317 VGND.n38 VGND.n12 0.1255
R318 VGND.n39 VGND.n11 0.1255
R319 VGND.n40 VGND.n10 0.1255
R320 VGND.n339 VGND.n48 0.1255
R321 VGND.n337 VGND.n50 0.1255
R322 VGND.n329 VGND.n58 0.1255
R323 VGND.n282 VGND.n230 0.124765
R324 VGND.n190 VGND.n128 0.124765
R325 VGND.n41 VGND.n9 0.124765
R326 VGND.n345 VGND.n344 0.124747
R327 VGND.n342 VGND.n45 0.124738
R328 VGND.n340 VGND.n47 0.124728
R329 VGND.n336 VGND.n51 0.124709
R330 VGND.n267 VGND.n246 0.124688
R331 VGND.n265 VGND.n248 0.124678
R332 VGND.n263 VGND.n250 0.124667
R333 VGND.n261 VGND.n252 0.124655
R334 VGND.n260 VGND.n253 0.124655
R335 VGND.n258 VGND.n255 0.124644
R336 VGND.n284 VGND.n228 0.124047
R337 VGND.n192 VGND.n126 0.124047
R338 VGND.n280 VGND.n232 0.124012
R339 VGND.n188 VGND.n130 0.124012
R340 VGND.n278 VGND.n234 0.123994
R341 VGND.n186 VGND.n132 0.123994
R342 VGND.n343 VGND.n6 0.123994
R343 VGND.n341 VGND.n46 0.123976
R344 VGND.n180 VGND.n138 0.123938
R345 VGND.n178 VGND.n140 0.123918
R346 VGND.n270 VGND.n243 0.123918
R347 VGND.n335 VGND.n52 0.123918
R348 VGND.n333 VGND.n54 0.123897
R349 VGND.n331 VGND.n56 0.123877
R350 VGND.n262 VGND.n251 0.123833
R351 VGND.n272 VGND.n271 0.123779
R352 VGND.n283 VGND.n229 0.12332
R353 VGND.n191 VGND.n127 0.12332
R354 VGND.n281 VGND.n231 0.123294
R355 VGND.n189 VGND.n129 0.123294
R356 VGND.n279 VGND.n233 0.123268
R357 VGND.n187 VGND.n131 0.123268
R358 VGND.n277 VGND.n235 0.123241
R359 VGND.n185 VGND.n133 0.123241
R360 VGND.n183 VGND.n135 0.123213
R361 VGND.n181 VGND.n137 0.123185
R362 VGND.n338 VGND.n49 0.123185
R363 VGND.n269 VGND.n244 0.123127
R364 VGND.n276 VGND.n236 0.122488
R365 VGND.n184 VGND.n134 0.122488
R366 VGND.n182 VGND.n136 0.122451
R367 VGND.n268 VGND.n245 0.122335
R368 VGND.n266 VGND.n247 0.122295
R369 VGND.n264 VGND.n249 0.122253
R370 VGND.n179 VGND.n139 0.121642
R371 VGND.n271 VGND.n242 0.121642
R372 VGND.n211 VGND.n210 0.120386
R373 VGND.n257 VGND.n94 0.115369
R374 VGND.n210 VGND.n209 0.112306
R375 VGND.n259 VGND.n258 0.111879
R376 VGND.n258 VGND.n257 0.111186
R377 VGND.n209 VGND.n208 0.109795
R378 VGND.n261 VGND.n260 0.108943
R379 VGND.n43 VGND.n42 0.108833
R380 VGND.n260 VGND.n259 0.107764
R381 VGND.n208 VGND.n207 0.107742
R382 VGND.n262 VGND.n261 0.107535
R383 VGND.n174 VGND.n140 0.107341
R384 VGND.n263 VGND.n262 0.106725
R385 VGND.n329 VGND.n328 0.106074
R386 VGND.n330 VGND.n329 0.105969
R387 VGND.n265 VGND.n264 0.1059
R388 VGND.n331 VGND.n330 0.105163
R389 VGND.n264 VGND.n263 0.104834
R390 VGND.n266 VGND.n265 0.104121
R391 VGND.n267 VGND.n266 0.103867
R392 VGND.n332 VGND.n331 0.10332
R393 VGND.n333 VGND.n332 0.10304
R394 VGND.n29 VGND.n28 0.102984
R395 VGND.n335 VGND.n334 0.102502
R396 VGND.n270 VGND.n269 0.102274
R397 VGND.n268 VGND.n267 0.10217
R398 VGND.n269 VGND.n268 0.101442
R399 VGND.n334 VGND.n333 0.101279
R400 VGND.n180 VGND.n179 0.1005
R401 VGND.n337 VGND.n336 0.100144
R402 VGND.n181 VGND.n180 0.0994435
R403 VGND.n338 VGND.n337 0.099433
R404 VGND.n336 VGND.n335 0.0992982
R405 VGND.n179 VGND.n178 0.0991552
R406 VGND.n271 VGND.n270 0.0991552
R407 VGND.n241 VGND.n238 0.0981562
R408 VGND.n275 VGND.n274 0.0977932
R409 VGND.n183 VGND.n182 0.0977932
R410 VGND.n340 VGND.n339 0.0976284
R411 VGND.n276 VGND.n275 0.0968228
R412 VGND.n184 VGND.n183 0.0968228
R413 VGND.n182 VGND.n181 0.0966929
R414 VGND.n341 VGND.n340 0.0965648
R415 VGND.n339 VGND.n338 0.0962384
R416 VGND.n277 VGND.n276 0.0962186
R417 VGND.n185 VGND.n184 0.0962186
R418 VGND.n254 VGND.n253 0.0959861
R419 VGND.n278 VGND.n277 0.0956231
R420 VGND.n186 VGND.n185 0.0956231
R421 VGND.n342 VGND.n341 0.0955348
R422 VGND.n343 VGND.n342 0.0948777
R423 VGND.n255 VGND.n254 0.0946781
R424 VGND.n31 VGND.n30 0.0945657
R425 VGND.n28 VGND.n27 0.0938949
R426 VGND.n206 VGND.n205 0.0937672
R427 VGND.n30 VGND.n29 0.0931452
R428 VGND.n204 VGND.n203 0.0930016
R429 VGND.n275 VGND.n237 0.0927256
R430 VGND.n279 VGND.n278 0.0927181
R431 VGND.n187 VGND.n186 0.0927181
R432 VGND.n207 VGND.n206 0.0923627
R433 VGND.n7 VGND.n5 0.0921667
R434 VGND.n280 VGND.n279 0.0920855
R435 VGND.n188 VGND.n187 0.0920855
R436 VGND.n344 VGND.n343 0.0919467
R437 VGND.n205 VGND.n204 0.0914722
R438 VGND.n344 VGND.n44 0.0912494
R439 VGND.n281 VGND.n280 0.091171
R440 VGND.n189 VGND.n188 0.091171
R441 VGND.n32 VGND.n31 0.0904148
R442 VGND.n252 VGND.n251 0.090027
R443 VGND.n253 VGND.n252 0.090027
R444 VGND.n282 VGND.n281 0.0898264
R445 VGND.n190 VGND.n189 0.0898264
R446 VGND.n284 VGND.n283 0.0891127
R447 VGND.n192 VGND.n191 0.0891127
R448 VGND.n38 VGND.n37 0.0881565
R449 VGND.n42 VGND.n41 0.0881488
R450 VGND.n41 VGND.n40 0.0879493
R451 VGND.n285 VGND.n284 0.0878131
R452 VGND.n193 VGND.n192 0.0878131
R453 VGND.n283 VGND.n282 0.0876124
R454 VGND.n191 VGND.n190 0.0876124
R455 VGND.n33 VGND.n32 0.0875536
R456 VGND.n251 VGND.n250 0.0871667
R457 VGND.n37 VGND.n36 0.0868953
R458 VGND.n326 VGND.n59 0.0866486
R459 VGND.n36 VGND.n35 0.0863769
R460 VGND.n202 VGND.n201 0.0859735
R461 VGND.n35 VGND.n34 0.0856762
R462 VGND.n44 VGND.n5 0.085541
R463 VGND.n250 VGND.n249 0.0855
R464 VGND.n34 VGND.n33 0.0852048
R465 VGND.n203 VGND.n202 0.0851591
R466 VGND.n40 VGND.n39 0.0850588
R467 VGND.n59 VGND.n58 0.0838333
R468 VGND.n292 VGND.n291 0.0835966
R469 VGND.n201 VGND.n200 0.0835966
R470 VGND.n288 VGND.n287 0.0833636
R471 VGND.n286 VGND.n285 0.0833488
R472 VGND.n194 VGND.n193 0.0833488
R473 VGND.n39 VGND.n38 0.0833488
R474 VGND.n289 VGND.n288 0.0825455
R475 VGND.n58 VGND.n57 0.0821667
R476 VGND.n196 VGND.n195 0.081981
R477 VGND.n290 VGND.n289 0.0819394
R478 VGND.n199 VGND.n198 0.0819394
R479 VGND.n287 VGND.n286 0.0816782
R480 VGND.n195 VGND.n194 0.0816782
R481 VGND.n249 VGND.n248 0.0816688
R482 VGND.n291 VGND.n290 0.0813424
R483 VGND.n200 VGND.n199 0.0813424
R484 VGND.n248 VGND.n247 0.0810921
R485 VGND.n272 VGND.n241 0.0797137
R486 VGND.n313 VGND.n94 0.0796453
R487 VGND.n256 VGND.n255 0.0796157
R488 VGND.n57 VGND.n56 0.0784221
R489 VGND.n56 VGND.n55 0.0778026
R490 VGND.n247 VGND.n246 0.0774231
R491 VGND.n246 VGND.n245 0.0767987
R492 VGND.n257 VGND.n256 0.0762042
R493 VGND.n55 VGND.n54 0.074218
R494 VGND.n54 VGND.n53 0.073552
R495 VGND.n245 VGND.n244 0.0732848
R496 VGND.n294 VGND.n220 0.0732142
R497 VGND.n292 VGND.n220 0.0719286
R498 VGND.n244 VGND.n243 0.0717025
R499 VGND.n140 VGND.n139 0.0701203
R500 VGND.n243 VGND.n242 0.0701203
R501 VGND.n53 VGND.n52 0.0701203
R502 VGND.n52 VGND.n51 0.068538
R503 VGND.n51 VGND.n50 0.0669557
R504 VGND.n139 VGND.n138 0.066858
R505 VGND.n242 VGND.n241 0.066858
R506 VGND.n237 VGND.n236 0.0667809
R507 VGND.n138 VGND.n137 0.066125
R508 VGND.n137 VGND.n136 0.0637716
R509 VGND.n50 VGND.n49 0.0637716
R510 VGND.n49 VGND.n48 0.063
R511 VGND.n136 VGND.n135 0.0614756
R512 VGND.n198 VGND.n197 0.0609482
R513 VGND.n48 VGND.n47 0.0606852
R514 VGND.n135 VGND.n134 0.0599512
R515 VGND.n47 VGND.n46 0.0584268
R516 VGND.n236 VGND.n235 0.0577289
R517 VGND.n134 VGND.n133 0.0577289
R518 VGND.n46 VGND.n45 0.0569024
R519 VGND.n235 VGND.n234 0.0562229
R520 VGND.n133 VGND.n132 0.0562229
R521 VGND.n219 VGND 0.0560556
R522 VGND.n122 VGND 0.0560556
R523 VGND.n172 VGND 0.0560556
R524 VGND.n161 VGND 0.0560556
R525 VGND.n176 VGND 0.0560556
R526 VGND.n297 VGND 0.0560556
R527 VGND.n240 VGND 0.0560556
R528 VGND.n312 VGND 0.0560556
R529 VGND.n316 VGND 0.0560556
R530 VGND.n90 VGND 0.0560556
R531 VGND.n314 VGND.n313 0.0554302
R532 VGND.n234 VGND.n233 0.0547169
R533 VGND.n132 VGND.n131 0.0547169
R534 VGND.n45 VGND.n6 0.0547169
R535 VGND.n345 VGND.n6 0.0532108
R536 VGND.n233 VGND.n232 0.0525833
R537 VGND.n131 VGND.n130 0.0525833
R538 VGND.n256 VGND.n93 0.0514752
R539 VGND.n232 VGND.n231 0.0510952
R540 VGND.n130 VGND.n129 0.0510952
R541 VGND.n231 VGND.n230 0.0490294
R542 VGND.n129 VGND.n128 0.0490294
R543 VGND.n294 VGND.n293 0.0488306
R544 VGND.n8 VGND.n7 0.046631
R545 VGND.n274 VGND.n238 0.0461288
R546 VGND.n230 VGND.n229 0.0460882
R547 VGND.n128 VGND.n127 0.0460882
R548 VGND.n9 VGND.n8 0.0460882
R549 VGND.n229 VGND.n228 0.0455581
R550 VGND.n127 VGND.n126 0.0455581
R551 VGND.n10 VGND.n9 0.0446176
R552 VGND.n228 VGND.n227 0.0441047
R553 VGND.n126 VGND.n125 0.0441047
R554 VGND.n227 VGND.n226 0.0411977
R555 VGND.n226 VGND.n225 0.0411977
R556 VGND.n125 VGND.n124 0.0411977
R557 VGND.n124 VGND.n123 0.0411977
R558 VGND.n12 VGND.n11 0.0411977
R559 VGND.n11 VGND.n10 0.0411977
R560 VGND.n327 VGND.n326 0.0401474
R561 VGND.n13 VGND.n12 0.0382907
R562 VGND.n94 VGND.n93 0.0381773
R563 VGND.n225 VGND.n224 0.0378563
R564 VGND.n123 VGND.n119 0.0378563
R565 VGND.n14 VGND.n13 0.0368372
R566 VGND.n224 VGND.n223 0.0364195
R567 VGND.n119 VGND.n118 0.0364195
R568 VGND.n345 VGND.n5 0.0353361
R569 VGND.n178 VGND.n177 0.0353101
R570 VGND.n15 VGND.n14 0.0349828
R571 VGND.n223 VGND.n222 0.0345909
R572 VGND.n118 VGND.n117 0.0345909
R573 VGND.n16 VGND.n15 0.033546
R574 VGND.n222 VGND.n221 0.0331705
R575 VGND.n117 VGND.n116 0.0331705
R576 VGND.n293 VGND.n221 0.03175
R577 VGND.n116 VGND.n115 0.03175
R578 VGND.n17 VGND.n16 0.03175
R579 VGND.n238 VGND.n237 0.0315583
R580 VGND.n115 VGND.n114 0.0303295
R581 VGND.n18 VGND.n17 0.0303295
R582 VGND.n19 VGND.n18 0.0289091
R583 VGND.n114 VGND.n113 0.0285899
R584 VGND.n113 VGND.n112 0.0260682
R585 VGND.n20 VGND.n19 0.0260682
R586 VGND.n112 VGND.n111 0.0257809
R587 VGND.n21 VGND.n20 0.0257809
R588 VGND.n22 VGND.n21 0.0232273
R589 VGND.n110 VGND.n109 0.0229719
R590 VGND.n23 VGND.n22 0.0229719
R591 VGND.n111 VGND.n110 0.0227222
R592 VGND.n109 VGND.n108 0.0201629
R593 VGND.n25 VGND.n23 0.0199444
R594 VGND.n108 VGND.n107 0.0185556
R595 VGND.n107 VGND.n106 0.0171667
R596 VGND.n92 VGND.n91 0.0169225
R597 VGND.n274 VGND.n273 0.0158374
R598 VGND.n106 VGND.n105 0.0157778
R599 VGND.n105 VGND.n104 0.013
R600 VGND.n104 VGND.n103 0.013
R601 VGND.n103 VGND.n102 0.0102222
R602 VGND.n26 VGND.n25 0.00911038
R603 VGND.n216 VGND.n102 0.00874176
R604 VGND.n295 VGND.n217 0.00816087
R605 VGND.n217 VGND.n216 0.00744444
R606 VGND.n197 VGND.n196 0.00285443
R607 VPWR.n4 VPWR.t27 739.681
R608 VPWR.n229 VPWR.t37 739.681
R609 VPWR.n231 VPWR.t11 739.681
R610 VPWR.n140 VPWR.t39 739.681
R611 VPWR.n138 VPWR.t1 739.681
R612 VPWR.n87 VPWR.t41 739.681
R613 VPWR.n8 VPWR.t33 739.681
R614 VPWR.n88 VPWR.t31 739.681
R615 VPWR.n112 VPWR.t29 739.681
R616 VPWR.n1 VPWR.t19 739.681
R617 VPWR.n0 VPWR.t15 739.681
R618 VPWR.n143 VPWR.t23 739.681
R619 VPWR.n85 VPWR.t13 739.681
R620 VPWR.n83 VPWR.t3 739.681
R621 VPWR.n56 VPWR.t35 739.681
R622 VPWR.n33 VPWR.t7 739.681
R623 VPWR.n12 VPWR.t9 739.681
R624 VPWR.n9 VPWR.t5 739.681
R625 VPWR.n6 VPWR.t17 739.681
R626 VPWR.n59 VPWR.t21 739.681
R627 VPWR.n149 VPWR.t25 739.681
R628 VPWR.n4 VPWR.t26 707.852
R629 VPWR.n229 VPWR.t36 707.852
R630 VPWR.n231 VPWR.t10 707.852
R631 VPWR.n140 VPWR.t38 707.852
R632 VPWR.n138 VPWR.t0 707.852
R633 VPWR.n143 VPWR.t22 707.852
R634 VPWR.n87 VPWR.t40 707.852
R635 VPWR.n85 VPWR.t12 707.852
R636 VPWR.n83 VPWR.t2 707.852
R637 VPWR.n56 VPWR.t34 707.852
R638 VPWR.n33 VPWR.t6 707.852
R639 VPWR.n12 VPWR.t8 707.852
R640 VPWR.n9 VPWR.t4 707.852
R641 VPWR.n8 VPWR.t32 707.852
R642 VPWR.n6 VPWR.t16 707.852
R643 VPWR.n59 VPWR.t20 707.852
R644 VPWR.n149 VPWR.t24 707.852
R645 VPWR.n88 VPWR.t30 707.852
R646 VPWR.n112 VPWR.t28 707.852
R647 VPWR.n1 VPWR.t18 707.852
R648 VPWR.n0 VPWR.t14 707.852
R649 VPWR.n144 VPWR.n143 13.377
R650 VPWR.n86 VPWR.n85 13.377
R651 VPWR.n84 VPWR.n83 13.377
R652 VPWR.n57 VPWR.n56 13.377
R653 VPWR.n34 VPWR.n33 13.377
R654 VPWR.n13 VPWR.n12 13.377
R655 VPWR.n10 VPWR.n9 13.377
R656 VPWR.n7 VPWR.n6 13.377
R657 VPWR.n60 VPWR.n59 13.377
R658 VPWR.n150 VPWR.n149 13.377
R659 VPWR VPWR.n4 13.3202
R660 VPWR.n230 VPWR.n229 13.3202
R661 VPWR VPWR.n231 13.3202
R662 VPWR VPWR.n140 13.3202
R663 VPWR.n139 VPWR.n138 13.3202
R664 VPWR VPWR.n87 13.3202
R665 VPWR VPWR.n8 13.3202
R666 VPWR.n89 VPWR.n88 13.3202
R667 VPWR.n113 VPWR.n112 13.3202
R668 VPWR.n2 VPWR.n1 13.3202
R669 VPWR.n235 VPWR.n0 13.3202
R670 VPWR.n228 VPWR 9.7375
R671 VPWR.n232 VPWR 9.39357
R672 VPWR.n145 VPWR.n144 8.51977
R673 VPWR.n222 VPWR 8.13646
R674 VPWR.n234 VPWR.n233 7.53241
R675 VPWR.n147 VPWR.n86 7.53109
R676 VPWR.n148 VPWR.n84 7.45619
R677 VPWR.n141 VPWR 7.19357
R678 VPWR.n151 VPWR.n150 6.79323
R679 VPWR.n223 VPWR.n7 6.76538
R680 VPWR.n146 VPWR 6.40107
R681 VPWR.n235 VPWR.n234 6.34337
R682 VPWR.n3 VPWR.n2 6.19552
R683 VPWR.n232 VPWR.n230 6.1805
R684 VPWR.n221 VPWR.n10 6.08268
R685 VPWR.n233 VPWR.n228 6.07746
R686 VPWR.n61 VPWR.n60 6.01772
R687 VPWR.n219 VPWR.n13 6.01019
R688 VPWR.n35 VPWR.n34 5.71852
R689 VPWR.n58 VPWR.n57 5.65925
R690 VPWR.n114 VPWR.n113 5.44488
R691 VPWR.n90 VPWR.n89 5.3655
R692 VPWR.n141 VPWR.n139 5.233
R693 VPWR.n225 VPWR 5.15791
R694 VPWR.n221 VPWR.n220 4.17361
R695 VPWR.n145 VPWR.n142 4.09662
R696 VPWR.n176 VPWR.n175 3.07281
R697 VPWR.n233 VPWR.n232 1.25038
R698 VPWR.n142 VPWR.n137 1.04638
R699 VPWR.n146 VPWR.n145 0.926193
R700 VPWR.n234 VPWR.n3 0.897709
R701 VPWR.n147 VPWR.n146 0.877511
R702 VPWR.n214 VPWR.n213 0.861295
R703 VPWR.n222 VPWR.n221 0.838747
R704 VPWR.n223 VPWR.n222 0.810795
R705 VPWR.n228 VPWR.n227 0.786394
R706 VPWR.n152 VPWR.n148 0.69817
R707 VPWR.n115 VPWR.n3 0.574375
R708 VPWR.n148 VPWR.n147 0.53698
R709 VPWR.n215 VPWR.n214 0.507602
R710 VPWR.n175 VPWR.n174 0.491158
R711 VPWR.n142 VPWR.n141 0.456575
R712 VPWR.n216 VPWR.n215 0.391496
R713 VPWR.n177 VPWR.n176 0.380996
R714 VPWR.n224 VPWR.n5 0.341219
R715 VPWR.n216 VPWR.n11 0.325974
R716 VPWR.n115 VPWR.n114 0.323617
R717 VPWR.n220 VPWR.n11 0.320751
R718 VPWR.n178 VPWR.n177 0.263105
R719 VPWR.n179 VPWR.n178 0.23221
R720 VPWR.n218 VPWR.n11 0.198913
R721 VPWR.n217 VPWR.n216 0.195812
R722 VPWR.n180 VPWR.n179 0.193814
R723 VPWR.n215 VPWR.n14 0.192808
R724 VPWR.n214 VPWR.n15 0.189894
R725 VPWR.n227 VPWR.n5 0.188146
R726 VPWR.n181 VPWR.n180 0.183989
R727 VPWR.n153 VPWR.n152 0.169675
R728 VPWR.n174 VPWR.n173 0.168706
R729 VPWR.n176 VPWR.n55 0.162658
R730 VPWR.n182 VPWR.n181 0.157627
R731 VPWR.n17 VPWR.n16 0.154418
R732 VPWR.n151 VPWR.n82 0.154418
R733 VPWR.n198 VPWR.n31 0.153485
R734 VPWR.n183 VPWR.n182 0.148565
R735 VPWR.n92 VPWR.n91 0.147626
R736 VPWR.n177 VPWR.n54 0.143882
R737 VPWR.n178 VPWR.n53 0.142412
R738 VPWR.n180 VPWR.n51 0.140206
R739 VPWR.n179 VPWR.n52 0.140035
R740 VPWR.n182 VPWR.n49 0.139637
R741 VPWR.n181 VPWR.n50 0.139471
R742 VPWR.n117 VPWR.n110 0.137548
R743 VPWR.n184 VPWR.n47 0.137405
R744 VPWR.n183 VPWR.n48 0.137265
R745 VPWR.n119 VPWR.n108 0.136933
R746 VPWR.n185 VPWR.n46 0.136661
R747 VPWR.n116 VPWR.n111 0.136661
R748 VPWR.n211 VPWR.n18 0.136529
R749 VPWR.n154 VPWR.n81 0.136529
R750 VPWR.n118 VPWR.n109 0.136042
R751 VPWR.n186 VPWR.n45 0.135917
R752 VPWR.n184 VPWR.n183 0.135794
R753 VPWR.n172 VPWR.n63 0.135785
R754 VPWR.n134 VPWR.n93 0.135774
R755 VPWR.n123 VPWR.n104 0.135656
R756 VPWR.n212 VPWR.n17 0.13561
R757 VPWR.n153 VPWR.n82 0.13561
R758 VPWR.n122 VPWR.n105 0.135531
R759 VPWR.n120 VPWR.n107 0.135409
R760 VPWR.n130 VPWR.n97 0.135368
R761 VPWR.n209 VPWR.n20 0.135321
R762 VPWR.n156 VPWR.n79 0.135321
R763 VPWR.n188 VPWR.n43 0.135289
R764 VPWR.n128 VPWR.n99 0.13524
R765 VPWR.n125 VPWR.n102 0.134994
R766 VPWR.n135 VPWR.n92 0.134918
R767 VPWR.n132 VPWR.n95 0.134667
R768 VPWR.n187 VPWR.n44 0.134429
R769 VPWR.n126 VPWR.n101 0.134203
R770 VPWR.n191 VPWR.n40 0.133884
R771 VPWR.n190 VPWR.n41 0.133884
R772 VPWR.n121 VPWR.n106 0.133884
R773 VPWR.n189 VPWR.n42 0.133783
R774 VPWR.n199 VPWR.n30 0.133617
R775 VPWR.n166 VPWR.n69 0.133617
R776 VPWR.n210 VPWR.n19 0.133536
R777 VPWR.n155 VPWR.n80 0.133536
R778 VPWR.n207 VPWR.n22 0.133312
R779 VPWR.n194 VPWR.n37 0.133312
R780 VPWR.n171 VPWR.n64 0.133312
R781 VPWR.n158 VPWR.n77 0.133312
R782 VPWR.n205 VPWR.n24 0.133205
R783 VPWR.n161 VPWR.n74 0.133101
R784 VPWR.n133 VPWR.n94 0.133
R785 VPWR.n201 VPWR.n28 0.132901
R786 VPWR.n164 VPWR.n71 0.132901
R787 VPWR.n131 VPWR.n96 0.132901
R788 VPWR.n196 VPWR.n35 0.13262
R789 VPWR.n169 VPWR.n66 0.13262
R790 VPWR.n127 VPWR.n100 0.13262
R791 VPWR.n193 VPWR.n38 0.132444
R792 VPWR.n124 VPWR.n103 0.132444
R793 VPWR.n192 VPWR.n39 0.13236
R794 VPWR.n206 VPWR.n23 0.132349
R795 VPWR.n159 VPWR.n76 0.132349
R796 VPWR.n203 VPWR.n26 0.132167
R797 VPWR.n162 VPWR.n73 0.132167
R798 VPWR.n129 VPWR.n98 0.13191
R799 VPWR.n168 VPWR.n67 0.131829
R800 VPWR.n111 VPWR.n110 0.131701
R801 VPWR.n208 VPWR.n21 0.131576
R802 VPWR.n157 VPWR.n78 0.131576
R803 VPWR.n160 VPWR.n75 0.131412
R804 VPWR.n204 VPWR.n25 0.131333
R805 VPWR.n202 VPWR.n27 0.131257
R806 VPWR.n163 VPWR.n72 0.131257
R807 VPWR.n195 VPWR.n36 0.130901
R808 VPWR.n170 VPWR.n65 0.130901
R809 VPWR.n137 VPWR.n136 0.130756
R810 VPWR.n167 VPWR.n68 0.130247
R811 VPWR.n110 VPWR.n109 0.130144
R812 VPWR.n185 VPWR.n184 0.130052
R813 VPWR.n200 VPWR.n29 0.129506
R814 VPWR.n165 VPWR.n70 0.129506
R815 VPWR.n173 VPWR.n62 0.12922
R816 VPWR.n212 VPWR.n211 0.124945
R817 VPWR.n154 VPWR.n153 0.124945
R818 VPWR.n186 VPWR.n185 0.12426
R819 VPWR.n211 VPWR.n210 0.122959
R820 VPWR.n155 VPWR.n154 0.122959
R821 VPWR.n109 VPWR.n108 0.122756
R822 VPWR.n108 VPWR.n107 0.122197
R823 VPWR.n198 VPWR.n197 0.121074
R824 VPWR.n210 VPWR.n209 0.12023
R825 VPWR.n156 VPWR.n155 0.12023
R826 VPWR.n209 VPWR.n208 0.119565
R827 VPWR.n157 VPWR.n156 0.119565
R828 VPWR.n218 VPWR.n217 0.118556
R829 VPWR.n137 VPWR.n90 0.118474
R830 VPWR.n107 VPWR.n106 0.117381
R831 VPWR.n187 VPWR.n186 0.117018
R832 VPWR.n188 VPWR.n187 0.116571
R833 VPWR.n208 VPWR.n207 0.115278
R834 VPWR.n158 VPWR.n157 0.115278
R835 VPWR.n217 VPWR.n14 0.114758
R836 VPWR.n93 VPWR.n92 0.114696
R837 VPWR.n197 VPWR.n32 0.114511
R838 VPWR.n207 VPWR.n206 0.114352
R839 VPWR.n159 VPWR.n158 0.114352
R840 VPWR.n105 VPWR.n104 0.114094
R841 VPWR.n206 VPWR.n205 0.113756
R842 VPWR.n160 VPWR.n159 0.113235
R843 VPWR.n95 VPWR.n94 0.113192
R844 VPWR.n104 VPWR.n103 0.113154
R845 VPWR.n94 VPWR.n93 0.112678
R846 VPWR.n97 VPWR.n96 0.112433
R847 VPWR.n199 VPWR.n198 0.112207
R848 VPWR.n189 VPWR.n188 0.111422
R849 VPWR.n205 VPWR.n204 0.111333
R850 VPWR.n101 VPWR.n100 0.111285
R851 VPWR.n204 VPWR.n203 0.111081
R852 VPWR.n162 VPWR.n161 0.111081
R853 VPWR.n15 VPWR.n14 0.111077
R854 VPWR.n161 VPWR.n160 0.110429
R855 VPWR.n99 VPWR.n98 0.110229
R856 VPWR.n163 VPWR.n162 0.11011
R857 VPWR.n96 VPWR.n95 0.109923
R858 VPWR.n106 VPWR.n105 0.10979
R859 VPWR.n191 VPWR.n190 0.109555
R860 VPWR.n173 VPWR.n172 0.108951
R861 VPWR.n201 VPWR.n200 0.108673
R862 VPWR.n165 VPWR.n164 0.108673
R863 VPWR.n203 VPWR.n202 0.108622
R864 VPWR.n102 VPWR.n101 0.108359
R865 VPWR.n103 VPWR.n102 0.108286
R866 VPWR.n98 VPWR.n97 0.10823
R867 VPWR.n190 VPWR.n189 0.107819
R868 VPWR.n100 VPWR.n99 0.107643
R869 VPWR.n225 VPWR.n5 0.107643
R870 VPWR.n202 VPWR.n201 0.107267
R871 VPWR.n164 VPWR.n163 0.107267
R872 VPWR.n167 VPWR.n166 0.107106
R873 VPWR.n16 VPWR.n15 0.106561
R874 VPWR.n192 VPWR.n191 0.105203
R875 VPWR.n193 VPWR.n192 0.105131
R876 VPWR.n172 VPWR.n171 0.104693
R877 VPWR.n195 VPWR.n194 0.104583
R878 VPWR.n171 VPWR.n170 0.104583
R879 VPWR.n194 VPWR.n193 0.104127
R880 VPWR.n196 VPWR.n195 0.103965
R881 VPWR.n170 VPWR.n169 0.103965
R882 VPWR.n197 VPWR.n196 0.103813
R883 VPWR.n169 VPWR.n168 0.103813
R884 VPWR.n168 VPWR.n167 0.103788
R885 VPWR.n200 VPWR.n199 0.103439
R886 VPWR.n166 VPWR.n165 0.103439
R887 VPWR.n213 VPWR.n212 0.100519
R888 VPWR.n18 VPWR.n17 0.0979265
R889 VPWR.n82 VPWR.n81 0.0979265
R890 VPWR.n19 VPWR.n18 0.0960882
R891 VPWR.n81 VPWR.n80 0.0960882
R892 VPWR.n20 VPWR.n19 0.0915714
R893 VPWR.n80 VPWR.n79 0.0915714
R894 VPWR.n21 VPWR.n20 0.088
R895 VPWR.n79 VPWR.n78 0.088
R896 VPWR.n22 VPWR.n21 0.0855694
R897 VPWR.n78 VPWR.n77 0.0855694
R898 VPWR.n136 VPWR.n91 0.0849982
R899 VPWR.n213 VPWR.n16 0.0844552
R900 VPWR.n220 VPWR.n219 0.0832089
R901 VPWR.n23 VPWR.n22 0.0820972
R902 VPWR.n77 VPWR.n76 0.0820972
R903 VPWR.n24 VPWR.n23 0.0792671
R904 VPWR.n76 VPWR.n75 0.0792671
R905 VPWR.n25 VPWR.n24 0.0775548
R906 VPWR.n75 VPWR.n74 0.0765135
R907 VPWR.n136 VPWR.n135 0.0741301
R908 VPWR.n74 VPWR.n73 0.0731351
R909 VPWR.n135 VPWR.n134 0.0724178
R910 VPWR.n26 VPWR.n25 0.0721667
R911 VPWR.n27 VPWR.n26 0.0705
R912 VPWR.n73 VPWR.n72 0.0705
R913 VPWR.n134 VPWR.n133 0.0688333
R914 VPWR.n28 VPWR.n27 0.0679342
R915 VPWR.n72 VPWR.n71 0.0679342
R916 VPWR.n32 VPWR.n31 0.0676642
R917 VPWR.n133 VPWR.n132 0.0655
R918 VPWR.n29 VPWR.n28 0.0646447
R919 VPWR.n71 VPWR.n70 0.0646447
R920 VPWR.n132 VPWR.n131 0.0646447
R921 VPWR.n30 VPWR.n29 0.063
R922 VPWR.n70 VPWR.n69 0.063
R923 VPWR.n131 VPWR.n130 0.0597105
R924 VPWR.n31 VPWR.n30 0.0589416
R925 VPWR.n69 VPWR.n68 0.0589416
R926 VPWR.n130 VPWR.n129 0.0581923
R927 VPWR.n68 VPWR.n67 0.057462
R928 VPWR.n144 VPWR 0.0573182
R929 VPWR.n86 VPWR 0.0573182
R930 VPWR.n84 VPWR 0.0573182
R931 VPWR.n57 VPWR 0.0573182
R932 VPWR.n34 VPWR 0.0573182
R933 VPWR.n13 VPWR 0.0573182
R934 VPWR.n10 VPWR 0.0573182
R935 VPWR.n7 VPWR 0.0573182
R936 VPWR.n60 VPWR 0.0573182
R937 VPWR.n150 VPWR 0.0573182
R938 VPWR.n129 VPWR.n128 0.0556948
R939 VPWR.n67 VPWR.n66 0.0542975
R940 VPWR.n36 VPWR.n35 0.0527152
R941 VPWR.n66 VPWR.n65 0.0527152
R942 VPWR.n128 VPWR.n127 0.0527152
R943 VPWR.n230 VPWR 0.0505
R944 VPWR.n139 VPWR 0.0505
R945 VPWR.n89 VPWR 0.0505
R946 VPWR.n113 VPWR 0.0505
R947 VPWR.n2 VPWR 0.0505
R948 VPWR VPWR.n235 0.0505
R949 VPWR.n127 VPWR.n126 0.0495506
R950 VPWR.n37 VPWR.n36 0.0483395
R951 VPWR.n65 VPWR.n64 0.0483395
R952 VPWR.n126 VPWR.n125 0.0479684
R953 VPWR.n38 VPWR.n37 0.047375
R954 VPWR.n64 VPWR.n63 0.047375
R955 VPWR.n35 VPWR.n32 0.0472033
R956 VPWR.n63 VPWR.n62 0.0463861
R957 VPWR.n39 VPWR.n38 0.0452531
R958 VPWR.n125 VPWR.n124 0.0452531
R959 VPWR.n124 VPWR.n123 0.0426875
R960 VPWR.n40 VPWR.n39 0.0416585
R961 VPWR.n62 VPWR.n61 0.0406786
R962 VPWR.n91 VPWR.n90 0.039507
R963 VPWR.n123 VPWR.n122 0.0390802
R964 VPWR.n41 VPWR.n40 0.0386098
R965 VPWR.n42 VPWR.n41 0.0386098
R966 VPWR.n122 VPWR.n121 0.0386098
R967 VPWR.n121 VPWR.n120 0.035561
R968 VPWR.n43 VPWR.n42 0.0351386
R969 VPWR.n116 VPWR.n115 0.0350681
R970 VPWR.n120 VPWR.n119 0.0325122
R971 VPWR.n44 VPWR.n43 0.0321265
R972 VPWR.n119 VPWR.n118 0.0306205
R973 VPWR.n45 VPWR.n44 0.0302619
R974 VPWR.n118 VPWR.n117 0.0276084
R975 VPWR.n46 VPWR.n45 0.0272857
R976 VPWR.n47 VPWR.n46 0.0257976
R977 VPWR.n117 VPWR.n116 0.0257976
R978 VPWR.n58 VPWR.n55 0.0244583
R979 VPWR.n48 VPWR.n47 0.0243095
R980 VPWR.n226 VPWR.n225 0.0243095
R981 VPWR.n175 VPWR.n58 0.0239375
R982 VPWR.n174 VPWR.n61 0.0227865
R983 VPWR.n227 VPWR.n226 0.0214028
R984 VPWR.n49 VPWR.n48 0.0210882
R985 VPWR.n50 VPWR.n49 0.0198452
R986 VPWR.n51 VPWR.n50 0.0166765
R987 VPWR.n52 VPWR.n51 0.0152059
R988 VPWR.n224 VPWR.n223 0.01479
R989 VPWR.n114 VPWR.n111 0.0131488
R990 VPWR.n226 VPWR.n224 0.0124293
R991 VPWR.n53 VPWR.n52 0.0121279
R992 VPWR.n54 VPWR.n53 0.0107941
R993 VPWR.n152 VPWR.n151 0.0104434
R994 VPWR.n55 VPWR.n54 0.00785294
R995 VPWR.n219 VPWR.n218 0.00590163
C0 uo_out[0] VGND 8.8973f
C1 VPWR VGND 0.149095p
C2 ring_0/skullfet_inverter_16.A VGND 4.53396f
C3 ring_0/skullfet_inverter_17.A VGND 4.70918f
C4 ring_0/skullfet_inverter_15.A VGND 4.82841f
C5 ring_0/skullfet_inverter_18.A VGND 4.90629f
C6 ring_0/skullfet_inverter_14.A VGND 4.98419f
C7 ring_0/skullfet_inverter_19.A VGND 4.923029f
C8 ring_0/skullfet_inverter_13.A VGND 4.78946f
C9 ring_0/skullfet_inverter_20.A VGND 4.72064f
C10 ring_0/skullfet_inverter_12.A VGND 5.60339f
C11 ring_0/skullfet_inverter_20.Y VGND 5.35745f
C12 ring_0/skullfet_inverter_11.A VGND 4.97718f
C13 ring_0/skullfet_inverter_1.A VGND 5.16765f
C14 ring_0/skullfet_inverter_10.A VGND 5.58737f
C15 ring_0/skullfet_inverter_2.A VGND 5.65285f
C16 ring_0/skullfet_inverter_9.A VGND 4.78733f
C17 ring_0/skullfet_inverter_3.A VGND 4.92041f
C18 ring_0/skullfet_inverter_4.A VGND 4.93544f
C19 ring_0/skullfet_inverter_8.A VGND 4.94116f
C20 ring_0/skullfet_inverter_7.A VGND 4.81796f
C21 ring_0/skullfet_inverter_6.A VGND 4.53217f
.ends

