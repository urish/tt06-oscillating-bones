magic
tech sky130A
magscale 1 2
timestamp 1712832449
<< viali >>
rect 5586 352 5620 386
rect 7519 352 7553 386
rect 9450 352 9484 386
rect 3934 263 3978 340
rect 4192 268 4226 302
rect 5866 263 5900 297
rect 6125 268 6159 302
rect 7798 263 7832 297
rect 8056 268 8090 302
rect 5299 153 5333 187
rect 7231 153 7265 187
rect 9146 132 9208 184
<< metal1 >>
rect 5574 386 5632 392
rect 5574 352 5586 386
rect 5620 352 5632 386
rect 3928 340 3984 352
rect 5574 346 5632 352
rect 7507 386 7565 392
rect 7507 352 7519 386
rect 7553 352 7565 386
rect 7507 346 7565 352
rect 9438 386 9496 392
rect 9438 352 9450 386
rect 9484 352 9496 386
rect 9438 346 9496 352
rect 3924 263 3934 340
rect 3986 263 3996 340
rect 4180 302 4238 308
rect 4180 268 4192 302
rect 4226 300 4238 302
rect 5582 300 5610 346
rect 4226 272 5610 300
rect 5854 297 5912 303
rect 4226 268 4238 272
rect 3928 251 3984 263
rect 4180 262 4238 268
rect 5854 263 5866 297
rect 5900 263 5912 297
rect 5854 257 5912 263
rect 6113 302 6171 308
rect 6113 268 6125 302
rect 6159 300 6171 302
rect 7515 300 7543 346
rect 6159 272 7543 300
rect 7786 297 7844 303
rect 6159 268 6171 272
rect 6113 262 6171 268
rect 7786 263 7798 297
rect 7832 263 7844 297
rect 7786 257 7844 263
rect 8044 302 8102 308
rect 8044 268 8056 302
rect 8090 300 8102 302
rect 9446 300 9474 346
rect 8090 272 9474 300
rect 8090 268 8102 272
rect 8044 262 8102 268
rect 5274 144 5284 196
rect 5346 187 5356 196
rect 5866 187 5900 257
rect 5346 153 5900 187
rect 7219 187 7277 193
rect 7798 187 7832 257
rect 7219 176 7231 187
rect 7265 176 7832 187
rect 5346 144 5356 153
rect 7202 124 7212 176
rect 7274 153 7832 176
rect 9134 184 9220 190
rect 7274 124 7284 153
rect 9134 132 9146 184
rect 9208 132 9220 184
rect 9134 126 9220 132
<< via1 >>
rect 3934 263 3978 340
rect 3978 263 3986 340
rect 5284 187 5346 196
rect 5284 153 5299 187
rect 5299 153 5333 187
rect 5333 153 5346 187
rect 5284 144 5346 153
rect 7212 153 7231 176
rect 7231 153 7265 176
rect 7265 153 7274 176
rect 7212 124 7274 153
rect 9146 132 9208 184
<< metal2 >>
rect 3920 340 4012 374
rect 3920 263 3934 340
rect 3986 263 4012 340
rect 3920 243 4012 263
rect 5284 196 5346 206
rect 5284 134 5346 144
rect 7212 176 7274 186
rect 7212 114 7274 124
rect 9146 184 9208 194
rect 9146 122 9208 132
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1701704242
transform 1 0 3902 0 1 48
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_2
timestamp 1701704242
transform 1 0 5834 0 1 48
box -38 -48 1786 592
use sky130_fd_sc_hd__dfxbp_1  sky130_fd_sc_hd__dfxbp_1_3
timestamp 1701704242
transform 1 0 7766 0 1 48
box -38 -48 1786 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1712785652
transform 1 0 5650 0 1 48
box -38 -48 222 592
use sky130_fd_sc_hd__tap_2  sky130_fd_sc_hd__tap_2_2
timestamp 1712785652
transform 1 0 7582 0 1 48
box -38 -48 222 592
<< labels >>
flabel metal2 3986 243 4012 374 1 FreeSans 2 0 0 0 IN
port 1 nsew default input
flabel metal2 5284 134 5346 206 1 FreeSans 2 0 0 0 ODIV2
port 2 nsew default output
flabel metal2 7212 114 7274 186 1 FreeSans 2 0 0 0 ODIV4
port 3 nsew default output
flabel metal2 9146 132 9208 184 1 FreeSans 2 0 0 0 ODIV8
port 4 nsew default output
<< end >>
