* NGSPICE file created from tt_um_oscillating_bones.ext - technology: sky130A

.subckt tt_um_oscillating_bones clk ena rst_n ui_in[0] ui_in[1] ui_in[2] ui_in[3]
+ ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4]
+ uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4]
+ uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4]
+ uio_out[5] uio_out[6] uio_out[7] uo_out[2] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VGND uo_out[0] uo_out[1] uo_out[3] VPWR
X0 a_13289_43697# uo_out[2].t2 VPWR.t47 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X1 a_16868_43697# a_17160_43997# a_17111_44089# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X2 a_16596_43697# a_16868_43697# VGND.t60 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X3 VPWR.t16 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X4 VGND.t7 uo_out[0].t2 ring_0/skullfet_inverter_6.A VGND.t6 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X5 a_17360_43697# a_17160_43997# a_17509_43723# VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X6 VGND.t46 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X7 VGND.t26 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_13.A VGND.t25 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X8 a_15221_43697# uo_out[1].t2 VPWR.t8 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X9 VPWR.t18 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X10 a_15179_44089# a_14664_43697# VPWR.t68 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X11 VGND.t76 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_20.A VGND.t75 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X12 ring_0/skullfet_inverter_6.A uo_out[0].t3 VPWR.t7 VPWR.t6 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X13 a_15577_43723# a_15357_43723# VGND.t82 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X14 VGND.t79 a_14664_43697# uo_out[2].t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X15 VPWR.t46 a_13289_43697# a_13296_43997# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X16 VGND.t61 a_15221_43697# a_15228_43997# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X17 VGND.t52 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_3.A VGND.t51 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X18 a_13843_43723# a_13296_43997# a_13496_43697# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X19 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_12.A VPWR.t22 VPWR.t21 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X20 VGND.t42 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_8.A VGND.t41 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X21 a_16501_43697# a_16596_43697# VGND.t59 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X22 a_12637_43697# a_12732_43697# VPWR.t32 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X23 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_15.A VGND.t15 VGND.t14 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X24 VGND.t68 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_12.A VGND.t67 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X25 a_17289_43723# a_17153_43697# a_16868_43697# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X26 a_13224_43723# a_12732_43697# VGND.t40 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X27 VPWR.t67 a_14664_43697# uo_out[2].t1 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X28 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_14.A VGND.t28 VGND.t27 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X29 VPWR.t61 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_18.A VPWR.t60 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X30 VGND.t70 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_2.A VGND.t69 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X31 a_17707_43723# a_17153_43697# a_17360_43697# VGND.t66 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X32 VGND.t13 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_1.A VGND.t12 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X33 a_15156_43723# a_14664_43697# VGND.t78 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
X34 a_14936_43697# a_15228_43997# a_15179_44089# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X35 a_13289_43697# uo_out[2].t3 VGND.t54 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X36 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_7.A VPWR.t36 VPWR.t35 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X37 ring_0/skullfet_inverter_12.A ring_0/skullfet_inverter_11.A VPWR.t57 VPWR.t56 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X38 ring_0/skullfet_inverter_2.A ring_0/skullfet_inverter_1.A VPWR.t59 VPWR.t58 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X39 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_8.A VPWR.t38 VPWR.t37 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X40 VGND.t11 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X41 a_14664_43697# a_14936_43697# VGND.t1 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X42 a_15428_43697# a_15228_43997# a_15577_43723# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X43 VGND.t18 a_12637_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X44 VGND.t47 a_13496_43697# a_13425_43723# VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X45 a_13247_44089# a_12732_43697# VPWR.t34 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X46 a_15221_43697# uo_out[1].t3 VGND.t9 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X47 a_16868_43697# a_17153_43697# a_17088_43723# VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X48 a_13645_43723# a_13425_43723# VGND.t34 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X49 VPWR.t29 ring_0/skullfet_inverter_16.A ring_0/skullfet_inverter_17.A VPWR.t28 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X50 VPWR.t70 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_19.A VPWR.t69 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X51 VGND.t36 a_15428_43697# a_15357_43723# VGND.t35 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X52 VGND.t39 a_12732_43697# uo_out[3].t0 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X53 VGND.t17 ring_0/skullfet_inverter_6.A ring_0/skullfet_inverter_7.A VGND.t16 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X54 VPWR.t17 a_17360_43697# a_17289_43723# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X55 a_14664_43697# a_14936_43697# VPWR.t0 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X56 VGND.t53 a_13289_43697# a_13296_43997# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X57 ring_0/skullfet_inverter_1.A ring_0/skullfet_inverter_20.Y VPWR.t11 VPWR.t10 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X58 VPWR.t13 ring_0/skullfet_inverter_15.A ring_0/skullfet_inverter_16.A VPWR.t12 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X59 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_19.A VPWR.t65 VPWR.t64 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X60 a_14569_43697# a_14664_43697# VGND.t77 VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X61 a_15604_44089# a_15357_43723# VPWR.t71 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X62 a_15357_43723# a_15221_43697# a_14936_43697# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X63 a_15428_43697# a_15221_43697# a_15604_44089# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X64 a_12732_43697# a_13004_43697# VGND.t31 VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.169 pd=1.82 as=0.08775 ps=0.92 w=0.65 l=0.15
X65 VGND.t3 ring_0/skullfet_inverter_4.A uo_out[0].t0 VGND.t2 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X66 a_17289_43723# a_17160_43997# a_16868_43697# VGND.t65 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X67 VPWR.t9 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N a_17707_43723# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X68 VPWR.t33 a_12732_43697# uo_out[3].t1 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X69 VGND.t30 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_11.A VGND.t29 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X70 ring_0/skullfet_inverter_10.A ring_0/skullfet_inverter_9.A VPWR.t4 VPWR.t3 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X71 VPWR.t20 ring_0/skullfet_inverter_13.A ring_0/skullfet_inverter_14.A VPWR.t19 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X72 ring_0/skullfet_inverter_7.A ring_0/skullfet_inverter_6.A VPWR.t15 VPWR.t14 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X73 a_17153_43697# uo_out[0].t4 VPWR.t5 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.0864 ps=0.91 w=0.64 l=0.15
X74 a_17536_44089# a_17289_43723# VPWR.t54 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X75 a_15775_43723# a_15221_43697# a_15428_43697# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X76 a_17360_43697# a_17153_43697# a_17536_44089# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X77 a_17111_44089# a_16596_43697# VPWR.t50 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0882 pd=0.84 as=0.1113 ps=1.37 w=0.42 l=0.15
X78 a_13004_43697# a_13296_43997# a_13247_44089# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0567 pd=0.69 as=0.0882 ps=0.84 w=0.42 l=0.15
X79 VPWR.t43 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X80 a_12732_43697# a_13004_43697# VPWR.t27 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X81 VGND.t49 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_4.A VGND.t48 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X82 VGND.t62 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X83 a_13496_43697# a_13296_43997# a_13645_43723# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0621 pd=0.705 as=0.0696 ps=0.765 w=0.36 l=0.15
X84 uo_out[0].t1 ring_0/skullfet_inverter_4.A VPWR.t2 VPWR.t1 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X85 ring_0/skullfet_inverter_11.A ring_0/skullfet_inverter_10.A VPWR.t26 VPWR.t25 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X86 a_16501_43697# a_16596_43697# VPWR.t49 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X87 a_14936_43697# a_15221_43697# a_15156_43723# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X88 VPWR.t55 a_17153_43697# a_17160_43997# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X89 VPWR.t31 a_15428_43697# a_15357_43723# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X90 VGND.t5 ring_0/skullfet_inverter_9.A ring_0/skullfet_inverter_10.A VGND.t4 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X91 ring_0/skullfet_inverter_4.A ring_0/skullfet_inverter_3.A VPWR.t42 VPWR.t41 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X92 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_13.A VGND.t24 VGND.t23 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X93 a_13425_43723# a_13296_43997# a_13004_43697# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X94 ring_0/skullfet_inverter_20.Y ring_0/skullfet_inverter_20.A VPWR.t63 VPWR.t62 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X95 a_12637_43697# a_12732_43697# VGND.t38 VGND.t37 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.097 ps=0.975 w=0.42 l=0.15
X96 a_13672_44089# a_13425_43723# VPWR.t30 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.07665 pd=0.785 as=0.178875 ps=1.26 w=0.42 l=0.15
X97 ring_0/skullfet_inverter_18.A ring_0/skullfet_inverter_17.A VGND.t72 VGND.t71 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X98 a_13425_43723# a_13289_43697# a_13004_43697# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1095 pd=1.075 as=0.0567 ps=0.69 w=0.42 l=0.15
X99 a_13496_43697# a_13289_43697# a_13672_44089# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.06825 pd=0.745 as=0.07665 ps=0.785 w=0.42 l=0.15
X100 VPWR.t39 a_14569_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.154 pd=1.335 as=0.26 ps=2.52 w=1 l=0.15
X101 a_15357_43723# a_15228_43997# a_14936_43697# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0989 pd=0.995 as=0.0684 ps=0.74 w=0.36 l=0.15
X102 VPWR.t53 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_2.Q_N a_15775_43723# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1092 pd=1.36 as=0.05775 ps=0.695 w=0.42 l=0.15
X103 VPWR.t24 ring_0/skullfet_inverter_14.A ring_0/skullfet_inverter_15.A VPWR.t23 sky130_fd_pr__pfet_01v8 ad=4.4307 pd=10.9 as=6.2694 ps=26.64 w=4.05 l=0.4
X104 a_17153_43697# uo_out[0].t5 VGND.t21 VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0567 ps=0.69 w=0.42 l=0.15
X105 a_13843_43723# a_13289_43697# a_13496_43697# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0813 pd=0.83 as=0.0621 ps=0.705 w=0.36 l=0.15
X106 a_17509_43723# a_17289_43723# VGND.t63 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.0696 pd=0.765 as=0.12095 ps=1.085 w=0.42 l=0.15
X107 VGND.t58 a_16596_43697# uo_out[1].t0 VGND.t57 sky130_fd_pr__nfet_01v8 ad=0.08775 pd=0.92 as=0.169 ps=1.82 w=0.65 l=0.15
X108 a_13004_43697# a_13289_43697# a_13224_43723# VGND.t43 sky130_fd_pr__nfet_01v8 ad=0.0684 pd=0.74 as=0.066 ps=0.745 w=0.36 l=0.15
X109 VGND.t20 a_17360_43697# a_17289_43723# VGND.t19 sky130_fd_pr__nfet_01v8 ad=0.12095 pd=1.085 as=0.0989 ps=0.995 w=0.64 l=0.15
X110 VGND.t50 a_16501_43697# freq_divider_0.sky130_fd_sc_hd__dfxbp_1_1.Q_N VGND.t0 sky130_fd_pr__nfet_01v8 ad=0.097 pd=0.975 as=0.169 ps=1.82 w=0.65 l=0.15
X111 VPWR.t52 a_15221_43697# a_15228_43997# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.0864 pd=0.91 as=0.1664 ps=1.8 w=0.64 l=0.15
X112 VGND.t22 freq_divider_0.sky130_fd_sc_hd__dfxbp_1_3.Q_N a_13843_43723# VGND.t8 sky130_fd_pr__nfet_01v8 ad=0.1092 pd=1.36 as=0.0813 ps=0.83 w=0.42 l=0.15
X113 a_15775_43723# a_15228_43997# a_15428_43697# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X114 ring_0/skullfet_inverter_19.A ring_0/skullfet_inverter_18.A VGND.t81 VGND.t80 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X115 a_16596_43697# a_16868_43697# VPWR.t51 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.27 pd=2.54 as=0.135 ps=1.27 w=1 l=0.15
X116 a_14569_43697# a_14664_43697# VPWR.t66 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.1664 pd=1.8 as=0.154 ps=1.335 w=0.64 l=0.15
X117 VGND.t74 ring_0/skullfet_inverter_20.A ring_0/skullfet_inverter_20.Y VGND.t73 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X118 ring_0/skullfet_inverter_17.A ring_0/skullfet_inverter_16.A VGND.t33 VGND.t32 sky130_fd_pr__nfet_01v8 ad=6.4314 pd=26.72 as=4.2687 ps=10.82 w=4.05 l=0.4
X119 a_17707_43723# a_17160_43997# a_17360_43697# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.05775 pd=0.695 as=0.06825 ps=0.745 w=0.42 l=0.15
X120 VPWR.t48 a_16596_43697# uo_out[1].t1 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.135 pd=1.27 as=0.26 ps=2.52 w=1 l=0.15
X121 VGND.t45 ring_0/skullfet_inverter_8.A ring_0/skullfet_inverter_9.A VGND.t44 sky130_fd_pr__nfet_01v8 ad=4.2687 pd=10.82 as=6.4314 ps=26.72 w=4.05 l=0.4
X122 VPWR.t40 a_13496_43697# a_13425_43723# freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB sky130_fd_pr__pfet_01v8_hvt ad=0.178875 pd=1.26 as=0.1095 ps=1.075 w=0.75 l=0.15
X123 ring_0/skullfet_inverter_3.A ring_0/skullfet_inverter_2.A VPWR.t45 VPWR.t44 sky130_fd_pr__pfet_01v8 ad=6.2694 pd=26.64 as=4.4307 ps=10.9 w=4.05 l=0.4
X124 VGND.t64 a_17153_43697# a_17160_43997# VGND.t10 sky130_fd_pr__nfet_01v8 ad=0.0567 pd=0.69 as=0.1092 ps=1.36 w=0.42 l=0.15
X125 a_17088_43723# a_16596_43697# VGND.t56 VGND.t55 sky130_fd_pr__nfet_01v8 ad=0.066 pd=0.745 as=0.1092 ps=1.36 w=0.42 l=0.15
R0 uo_out[2].n2 uo_out[2].t1 313.104
R1 uo_out[2].n0 uo_out[2].t2 294.557
R2 uo_out[2].t0 uo_out[2].n2 265.769
R3 uo_out[2] uo_out[2].t0 262.318
R4 uo_out[2].n0 uo_out[2].t3 211.01
R5 uo_out[2].n1 uo_out[2].n0 152
R6 uo_out[2].n5 uo_out[2] 12.1482
R7 uo_out[2].n4 uo_out[2].n1 11.6311
R8 uo_out[2].n4 uo_out[2].n3 9.3005
R9 uo_out[2].n3 uo_out[2] 7.17626
R10 uo_out[2].n3 uo_out[2].n2 4.84898
R11 uo_out[2].n5 uo_out[2].n4 4.51042
R12 uo_out[2].n1 uo_out[2] 1.37896
R13 uo_out[2] uo_out[2].n5 0.0730806
R14 VPWR.n112 VPWR.t63 739.681
R15 VPWR.n114 VPWR.t70 739.681
R16 VPWR.n116 VPWR.t65 739.681
R17 VPWR.n150 VPWR.t22 739.681
R18 VPWR.n148 VPWR.t20 739.681
R19 VPWR.n84 VPWR.t26 739.681
R20 VPWR.n5 VPWR.t59 739.681
R21 VPWR.n85 VPWR.t24 739.681
R22 VPWR.n109 VPWR.t13 739.681
R23 VPWR.n122 VPWR.t29 739.681
R24 VPWR.n119 VPWR.t61 739.681
R25 VPWR.n153 VPWR.t57 739.681
R26 VPWR.n82 VPWR.t4 739.681
R27 VPWR.n80 VPWR.t38 739.681
R28 VPWR.n53 VPWR.t7 739.681
R29 VPWR.n30 VPWR.t2 739.681
R30 VPWR.n9 VPWR.t42 739.681
R31 VPWR.n6 VPWR.t45 739.681
R32 VPWR.n3 VPWR.t11 739.681
R33 VPWR.n56 VPWR.t15 739.681
R34 VPWR.n159 VPWR.t36 739.681
R35 VPWR.n112 VPWR.t62 707.852
R36 VPWR.n114 VPWR.t69 707.852
R37 VPWR.n116 VPWR.t64 707.852
R38 VPWR.n150 VPWR.t21 707.852
R39 VPWR.n148 VPWR.t19 707.852
R40 VPWR.n153 VPWR.t56 707.852
R41 VPWR.n84 VPWR.t25 707.852
R42 VPWR.n82 VPWR.t3 707.852
R43 VPWR.n80 VPWR.t37 707.852
R44 VPWR.n53 VPWR.t6 707.852
R45 VPWR.n30 VPWR.t1 707.852
R46 VPWR.n9 VPWR.t41 707.852
R47 VPWR.n6 VPWR.t44 707.852
R48 VPWR.n5 VPWR.t58 707.852
R49 VPWR.n3 VPWR.t10 707.852
R50 VPWR.n56 VPWR.t14 707.852
R51 VPWR.n159 VPWR.t35 707.852
R52 VPWR.n85 VPWR.t23 707.852
R53 VPWR.n109 VPWR.t12 707.852
R54 VPWR.n122 VPWR.t28 707.852
R55 VPWR.n119 VPWR.t60 707.852
R56 VPWR.n285 VPWR.t34 667.734
R57 VPWR.n320 VPWR.t68 667.734
R58 VPWR.n354 VPWR.t50 667.734
R59 VPWR.n299 VPWR.t18 666.677
R60 VPWR.n334 VPWR.t53 666.677
R61 VPWR.n238 VPWR.t9 666.677
R62 VPWR.n304 VPWR.n303 604.394
R63 VPWR.n251 VPWR.n250 604.394
R64 VPWR.n372 VPWR.n371 604.394
R65 VPWR.n273 VPWR.n272 333.348
R66 VPWR.n261 VPWR.n260 333.348
R67 VPWR.n352 VPWR.n246 333.348
R68 VPWR.n292 VPWR.n269 320.976
R69 VPWR.n327 VPWR.n255 320.976
R70 VPWR.n243 VPWR.n242 320.976
R71 VPWR.n276 VPWR.n275 240.522
R72 VPWR.n263 VPWR.n262 240.522
R73 VPWR.n346 VPWR.n345 240.522
R74 VPWR.n269 VPWR.t30 113.98
R75 VPWR.n255 VPWR.t71 113.98
R76 VPWR.n242 VPWR.t54 113.98
R77 VPWR.n275 VPWR.t32 61.9872
R78 VPWR.n262 VPWR.t66 61.9872
R79 VPWR.n345 VPWR.t49 61.9872
R80 VPWR.n303 VPWR.t47 41.5552
R81 VPWR.n303 VPWR.t46 41.5552
R82 VPWR.n250 VPWR.t8 41.5552
R83 VPWR.n250 VPWR.t52 41.5552
R84 VPWR.n371 VPWR.t5 41.5552
R85 VPWR.n371 VPWR.t55 41.5552
R86 VPWR.n269 VPWR.t40 35.4605
R87 VPWR.n255 VPWR.t31 35.4605
R88 VPWR.n242 VPWR.t17 35.4605
R89 VPWR.n281 VPWR.n280 34.6358
R90 VPWR.n280 VPWR.n279 34.6358
R91 VPWR.n298 VPWR.n297 34.6358
R92 VPWR.n297 VPWR.n267 34.6358
R93 VPWR.n293 VPWR.n267 34.6358
R94 VPWR.n291 VPWR.n290 34.6358
R95 VPWR.n290 VPWR.n270 34.6358
R96 VPWR.n286 VPWR.n270 34.6358
R97 VPWR.n310 VPWR.n309 34.6358
R98 VPWR.n309 VPWR.n264 34.6358
R99 VPWR.n305 VPWR.n264 34.6358
R100 VPWR.n316 VPWR.n315 34.6358
R101 VPWR.n315 VPWR.n314 34.6358
R102 VPWR.n333 VPWR.n253 34.6358
R103 VPWR.n329 VPWR.n253 34.6358
R104 VPWR.n329 VPWR.n328 34.6358
R105 VPWR.n326 VPWR.n256 34.6358
R106 VPWR.n322 VPWR.n256 34.6358
R107 VPWR.n322 VPWR.n321 34.6358
R108 VPWR.n344 VPWR.n249 34.6358
R109 VPWR.n340 VPWR.n249 34.6358
R110 VPWR.n340 VPWR.n339 34.6358
R111 VPWR.n351 VPWR.n247 34.6358
R112 VPWR.n347 VPWR.n247 34.6358
R113 VPWR.n366 VPWR.n365 34.6358
R114 VPWR.n365 VPWR.n364 34.6358
R115 VPWR.n364 VPWR.n240 34.6358
R116 VPWR.n360 VPWR.n359 34.6358
R117 VPWR.n359 VPWR.n358 34.6358
R118 VPWR.n358 VPWR.n244 34.6358
R119 VPWR.n284 VPWR.n273 32.0005
R120 VPWR.n261 VPWR.n258 32.0005
R121 VPWR.n353 VPWR.n352 32.0005
R122 VPWR.n373 VPWR.n372 30.7593
R123 VPWR.n285 VPWR.n284 30.4946
R124 VPWR.n320 VPWR.n258 30.4946
R125 VPWR.n354 VPWR.n353 30.4946
R126 VPWR.n275 VPWR.t16 30.1692
R127 VPWR.n262 VPWR.t39 30.1692
R128 VPWR.n345 VPWR.t43 30.1692
R129 VPWR.n299 VPWR.n298 27.4829
R130 VPWR.n310 VPWR.n263 27.4829
R131 VPWR.n334 VPWR.n333 27.4829
R132 VPWR.n346 VPWR.n344 27.4829
R133 VPWR.n366 VPWR.n238 27.4829
R134 VPWR.n272 VPWR.t27 26.5955
R135 VPWR.n272 VPWR.t33 26.5955
R136 VPWR.n260 VPWR.t0 26.5955
R137 VPWR.n260 VPWR.t67 26.5955
R138 VPWR.n246 VPWR.t51 26.5955
R139 VPWR.n246 VPWR.t48 26.5955
R140 VPWR.n279 VPWR.n276 25.6005
R141 VPWR.n314 VPWR.n263 25.6005
R142 VPWR.n347 VPWR.n346 25.6005
R143 VPWR.n304 VPWR.n265 22.9652
R144 VPWR.n335 VPWR.n251 22.9652
R145 VPWR.n372 VPWR.n370 22.9652
R146 VPWR.n299 VPWR.n265 21.8358
R147 VPWR.n335 VPWR.n334 21.8358
R148 VPWR.n370 VPWR.n238 21.8358
R149 VPWR.n373 VPWR.n237 21.795
R150 VPWR.n305 VPWR.n304 21.4593
R151 VPWR.n339 VPWR.n251 21.4593
R152 VPWR.n293 VPWR.n292 18.4476
R153 VPWR.n328 VPWR.n327 18.4476
R154 VPWR.n243 VPWR.n240 18.4476
R155 VPWR.n292 VPWR.n291 16.1887
R156 VPWR.n327 VPWR.n326 16.1887
R157 VPWR.n360 VPWR.n243 16.1887
R158 VPWR.n286 VPWR.n285 15.0593
R159 VPWR.n321 VPWR.n320 15.0593
R160 VPWR.n354 VPWR.n244 15.0593
R161 VPWR.n154 VPWR.n153 13.377
R162 VPWR.n83 VPWR.n82 13.377
R163 VPWR.n81 VPWR.n80 13.377
R164 VPWR.n54 VPWR.n53 13.377
R165 VPWR.n31 VPWR.n30 13.377
R166 VPWR.n10 VPWR.n9 13.377
R167 VPWR.n7 VPWR.n6 13.377
R168 VPWR.n4 VPWR.n3 13.377
R169 VPWR.n57 VPWR.n56 13.377
R170 VPWR.n160 VPWR.n159 13.377
R171 VPWR VPWR.n112 13.3202
R172 VPWR.n115 VPWR.n114 13.3202
R173 VPWR VPWR.n116 13.3202
R174 VPWR VPWR.n150 13.3202
R175 VPWR.n149 VPWR.n148 13.3202
R176 VPWR VPWR.n84 13.3202
R177 VPWR VPWR.n5 13.3202
R178 VPWR.n86 VPWR.n85 13.3202
R179 VPWR.n110 VPWR.n109 13.3202
R180 VPWR.n123 VPWR.n122 13.3202
R181 VPWR.n120 VPWR.n119 13.3202
R182 VPWR.n113 VPWR 9.7375
R183 VPWR.n117 VPWR 9.39357
R184 VPWR.n372 VPWR.n0 9.3005
R185 VPWR.n370 VPWR.n369 9.3005
R186 VPWR.n368 VPWR.n238 9.3005
R187 VPWR.n367 VPWR.n366 9.3005
R188 VPWR.n365 VPWR.n239 9.3005
R189 VPWR.n364 VPWR.n363 9.3005
R190 VPWR.n362 VPWR.n240 9.3005
R191 VPWR.n361 VPWR.n360 9.3005
R192 VPWR.n359 VPWR.n241 9.3005
R193 VPWR.n358 VPWR.n357 9.3005
R194 VPWR.n356 VPWR.n244 9.3005
R195 VPWR.n355 VPWR.n354 9.3005
R196 VPWR.n353 VPWR.n245 9.3005
R197 VPWR.n351 VPWR.n350 9.3005
R198 VPWR.n349 VPWR.n247 9.3005
R199 VPWR.n348 VPWR.n347 9.3005
R200 VPWR.n346 VPWR.n248 9.3005
R201 VPWR.n344 VPWR.n343 9.3005
R202 VPWR.n342 VPWR.n249 9.3005
R203 VPWR.n341 VPWR.n340 9.3005
R204 VPWR.n339 VPWR.n338 9.3005
R205 VPWR.n337 VPWR.n251 9.3005
R206 VPWR.n336 VPWR.n335 9.3005
R207 VPWR.n334 VPWR.n252 9.3005
R208 VPWR.n333 VPWR.n332 9.3005
R209 VPWR.n331 VPWR.n253 9.3005
R210 VPWR.n330 VPWR.n329 9.3005
R211 VPWR.n328 VPWR.n254 9.3005
R212 VPWR.n326 VPWR.n325 9.3005
R213 VPWR.n324 VPWR.n256 9.3005
R214 VPWR.n323 VPWR.n322 9.3005
R215 VPWR.n321 VPWR.n257 9.3005
R216 VPWR.n320 VPWR.n319 9.3005
R217 VPWR.n318 VPWR.n258 9.3005
R218 VPWR.n317 VPWR.n316 9.3005
R219 VPWR.n315 VPWR.n259 9.3005
R220 VPWR.n314 VPWR.n313 9.3005
R221 VPWR.n312 VPWR.n263 9.3005
R222 VPWR.n311 VPWR.n310 9.3005
R223 VPWR.n309 VPWR.n308 9.3005
R224 VPWR.n307 VPWR.n264 9.3005
R225 VPWR.n306 VPWR.n305 9.3005
R226 VPWR.n304 VPWR.n302 9.3005
R227 VPWR.n301 VPWR.n265 9.3005
R228 VPWR.n300 VPWR.n299 9.3005
R229 VPWR.n298 VPWR.n266 9.3005
R230 VPWR.n297 VPWR.n296 9.3005
R231 VPWR.n295 VPWR.n267 9.3005
R232 VPWR.n294 VPWR.n293 9.3005
R233 VPWR.n291 VPWR.n268 9.3005
R234 VPWR.n290 VPWR.n289 9.3005
R235 VPWR.n288 VPWR.n270 9.3005
R236 VPWR.n287 VPWR.n286 9.3005
R237 VPWR.n285 VPWR.n271 9.3005
R238 VPWR.n284 VPWR.n283 9.3005
R239 VPWR.n282 VPWR.n281 9.3005
R240 VPWR.n280 VPWR.n274 9.3005
R241 VPWR.n279 VPWR.n278 9.3005
R242 VPWR.n155 VPWR.n154 8.51977
R243 VPWR.n232 VPWR 8.13646
R244 VPWR.n121 VPWR.n118 7.53241
R245 VPWR.n157 VPWR.n83 7.53109
R246 VPWR.n158 VPWR.n81 7.45619
R247 VPWR.n277 VPWR.n276 7.4049
R248 VPWR.n151 VPWR 7.19357
R249 VPWR.n161 VPWR.n160 6.79323
R250 VPWR.n233 VPWR.n4 6.76538
R251 VPWR.n156 VPWR 6.40107
R252 VPWR.n121 VPWR.n120 6.34337
R253 VPWR.n124 VPWR.n123 6.19552
R254 VPWR.n117 VPWR.n115 6.1805
R255 VPWR.n231 VPWR.n7 6.08268
R256 VPWR.n118 VPWR.n113 6.07746
R257 VPWR.n58 VPWR.n57 6.01772
R258 VPWR.n229 VPWR.n10 6.01019
R259 VPWR.n32 VPWR.n31 5.71852
R260 VPWR.n55 VPWR.n54 5.65925
R261 VPWR.n111 VPWR.n110 5.44488
R262 VPWR.n87 VPWR.n86 5.3655
R263 VPWR.n151 VPWR.n149 5.233
R264 VPWR.n231 VPWR.n230 4.17361
R265 VPWR.n155 VPWR.n152 4.09662
R266 VPWR.n237 VPWR 3.1965
R267 VPWR.n186 VPWR.n185 3.07281
R268 VPWR.n281 VPWR.n273 2.63579
R269 VPWR.n316 VPWR.n261 2.63579
R270 VPWR.n352 VPWR.n351 2.63579
R271 VPWR.n237 VPWR.n236 1.96192
R272 VPWR.n118 VPWR.n117 1.25038
R273 VPWR.n152 VPWR.n147 1.04638
R274 VPWR.n156 VPWR.n155 0.926193
R275 VPWR.n124 VPWR.n121 0.897709
R276 VPWR.n157 VPWR.n156 0.877511
R277 VPWR.n224 VPWR.n223 0.861295
R278 VPWR.n232 VPWR.n231 0.838747
R279 VPWR.n233 VPWR.n232 0.810795
R280 VPWR.n113 VPWR.n2 0.786394
R281 VPWR.n162 VPWR.n158 0.69817
R282 VPWR.n125 VPWR.n124 0.574375
R283 VPWR.n158 VPWR.n157 0.53698
R284 VPWR.n225 VPWR.n224 0.507602
R285 VPWR.n185 VPWR.n184 0.491158
R286 VPWR.n152 VPWR.n151 0.456575
R287 VPWR.n226 VPWR.n225 0.391496
R288 VPWR.n187 VPWR.n186 0.380996
R289 VPWR.n235 VPWR.n234 0.341219
R290 VPWR.n226 VPWR.n8 0.325974
R291 VPWR.n125 VPWR.n111 0.323617
R292 VPWR.n230 VPWR.n8 0.320751
R293 VPWR.n188 VPWR.n187 0.263105
R294 VPWR.n189 VPWR.n188 0.23221
R295 VPWR.n228 VPWR.n8 0.198913
R296 VPWR.n227 VPWR.n226 0.195812
R297 VPWR.n190 VPWR.n189 0.193814
R298 VPWR.n225 VPWR.n11 0.192808
R299 VPWR.n224 VPWR.n12 0.189894
R300 VPWR.n235 VPWR.n2 0.188146
R301 VPWR.n191 VPWR.n190 0.183989
R302 VPWR.n163 VPWR.n162 0.169675
R303 VPWR.n184 VPWR.n183 0.168706
R304 VPWR.n186 VPWR.n52 0.162658
R305 VPWR.n192 VPWR.n191 0.157627
R306 VPWR.n277 VPWR 0.156264
R307 VPWR.n14 VPWR.n13 0.154418
R308 VPWR.n161 VPWR.n79 0.154418
R309 VPWR.n208 VPWR.n28 0.153485
R310 VPWR.n193 VPWR.n192 0.148565
R311 VPWR.n89 VPWR.n88 0.147626
R312 VPWR.n278 VPWR.n277 0.144904
R313 VPWR.n187 VPWR.n51 0.143882
R314 VPWR.n188 VPWR.n50 0.142412
R315 VPWR.n190 VPWR.n48 0.140206
R316 VPWR.n189 VPWR.n49 0.140035
R317 VPWR.n192 VPWR.n46 0.139637
R318 VPWR.n191 VPWR.n47 0.139471
R319 VPWR.n127 VPWR.n107 0.137548
R320 VPWR.n194 VPWR.n44 0.137405
R321 VPWR.n193 VPWR.n45 0.137265
R322 VPWR.n129 VPWR.n105 0.136933
R323 VPWR.n195 VPWR.n43 0.136661
R324 VPWR.n126 VPWR.n108 0.136661
R325 VPWR.n221 VPWR.n15 0.136529
R326 VPWR.n164 VPWR.n78 0.136529
R327 VPWR.n128 VPWR.n106 0.136042
R328 VPWR.n196 VPWR.n42 0.135917
R329 VPWR.n194 VPWR.n193 0.135794
R330 VPWR.n182 VPWR.n60 0.135785
R331 VPWR.n144 VPWR.n90 0.135774
R332 VPWR.n133 VPWR.n101 0.135656
R333 VPWR.n222 VPWR.n14 0.13561
R334 VPWR.n163 VPWR.n79 0.13561
R335 VPWR.n132 VPWR.n102 0.135531
R336 VPWR.n130 VPWR.n104 0.135409
R337 VPWR.n140 VPWR.n94 0.135368
R338 VPWR.n219 VPWR.n17 0.135321
R339 VPWR.n166 VPWR.n76 0.135321
R340 VPWR.n198 VPWR.n40 0.135289
R341 VPWR.n138 VPWR.n96 0.13524
R342 VPWR.n135 VPWR.n99 0.134994
R343 VPWR.n145 VPWR.n89 0.134918
R344 VPWR.n142 VPWR.n92 0.134667
R345 VPWR.n197 VPWR.n41 0.134429
R346 VPWR.n136 VPWR.n98 0.134203
R347 VPWR.n201 VPWR.n37 0.133884
R348 VPWR.n200 VPWR.n38 0.133884
R349 VPWR.n131 VPWR.n103 0.133884
R350 VPWR.n199 VPWR.n39 0.133783
R351 VPWR.n209 VPWR.n27 0.133617
R352 VPWR.n176 VPWR.n66 0.133617
R353 VPWR.n220 VPWR.n16 0.133536
R354 VPWR.n165 VPWR.n77 0.133536
R355 VPWR.n217 VPWR.n19 0.133312
R356 VPWR.n204 VPWR.n34 0.133312
R357 VPWR.n181 VPWR.n61 0.133312
R358 VPWR.n168 VPWR.n74 0.133312
R359 VPWR.n215 VPWR.n21 0.133205
R360 VPWR.n171 VPWR.n71 0.133101
R361 VPWR.n143 VPWR.n91 0.133
R362 VPWR.n211 VPWR.n25 0.132901
R363 VPWR.n174 VPWR.n68 0.132901
R364 VPWR.n141 VPWR.n93 0.132901
R365 VPWR.n206 VPWR.n32 0.13262
R366 VPWR.n179 VPWR.n63 0.13262
R367 VPWR.n137 VPWR.n97 0.13262
R368 VPWR.n203 VPWR.n35 0.132444
R369 VPWR.n134 VPWR.n100 0.132444
R370 VPWR.n202 VPWR.n36 0.13236
R371 VPWR.n216 VPWR.n20 0.132349
R372 VPWR.n169 VPWR.n73 0.132349
R373 VPWR.n213 VPWR.n23 0.132167
R374 VPWR.n172 VPWR.n70 0.132167
R375 VPWR.n139 VPWR.n95 0.13191
R376 VPWR.n178 VPWR.n64 0.131829
R377 VPWR.n108 VPWR.n107 0.131701
R378 VPWR.n218 VPWR.n18 0.131576
R379 VPWR.n167 VPWR.n75 0.131576
R380 VPWR.n170 VPWR.n72 0.131412
R381 VPWR.n214 VPWR.n22 0.131333
R382 VPWR.n212 VPWR.n24 0.131257
R383 VPWR.n173 VPWR.n69 0.131257
R384 VPWR.n205 VPWR.n33 0.130901
R385 VPWR.n180 VPWR.n62 0.130901
R386 VPWR.n147 VPWR.n146 0.130756
R387 VPWR.n177 VPWR.n65 0.130247
R388 VPWR.n107 VPWR.n106 0.130144
R389 VPWR.n195 VPWR.n194 0.130052
R390 VPWR.n210 VPWR.n26 0.129506
R391 VPWR.n175 VPWR.n67 0.129506
R392 VPWR.n183 VPWR.n59 0.12922
R393 VPWR.n222 VPWR.n221 0.124945
R394 VPWR.n164 VPWR.n163 0.124945
R395 VPWR.n196 VPWR.n195 0.12426
R396 VPWR.n221 VPWR.n220 0.122959
R397 VPWR.n165 VPWR.n164 0.122959
R398 VPWR.n106 VPWR.n105 0.122756
R399 VPWR.n105 VPWR.n104 0.122197
R400 VPWR.n208 VPWR.n207 0.121074
R401 VPWR.n369 VPWR.n0 0.120292
R402 VPWR.n369 VPWR.n368 0.120292
R403 VPWR.n368 VPWR.n367 0.120292
R404 VPWR.n367 VPWR.n239 0.120292
R405 VPWR.n363 VPWR.n239 0.120292
R406 VPWR.n363 VPWR.n362 0.120292
R407 VPWR.n362 VPWR.n361 0.120292
R408 VPWR.n361 VPWR.n241 0.120292
R409 VPWR.n357 VPWR.n241 0.120292
R410 VPWR.n357 VPWR.n356 0.120292
R411 VPWR.n356 VPWR.n355 0.120292
R412 VPWR.n355 VPWR.n245 0.120292
R413 VPWR.n350 VPWR.n245 0.120292
R414 VPWR.n350 VPWR.n349 0.120292
R415 VPWR.n349 VPWR.n348 0.120292
R416 VPWR.n348 VPWR.n248 0.120292
R417 VPWR.n343 VPWR.n248 0.120292
R418 VPWR.n337 VPWR.n336 0.120292
R419 VPWR.n336 VPWR.n252 0.120292
R420 VPWR.n332 VPWR.n252 0.120292
R421 VPWR.n332 VPWR.n331 0.120292
R422 VPWR.n331 VPWR.n330 0.120292
R423 VPWR.n330 VPWR.n254 0.120292
R424 VPWR.n325 VPWR.n254 0.120292
R425 VPWR.n325 VPWR.n324 0.120292
R426 VPWR.n324 VPWR.n323 0.120292
R427 VPWR.n323 VPWR.n257 0.120292
R428 VPWR.n319 VPWR.n257 0.120292
R429 VPWR.n319 VPWR.n318 0.120292
R430 VPWR.n318 VPWR.n317 0.120292
R431 VPWR.n317 VPWR.n259 0.120292
R432 VPWR.n313 VPWR.n259 0.120292
R433 VPWR.n313 VPWR.n312 0.120292
R434 VPWR.n312 VPWR.n311 0.120292
R435 VPWR.n302 VPWR.n301 0.120292
R436 VPWR.n301 VPWR.n300 0.120292
R437 VPWR.n300 VPWR.n266 0.120292
R438 VPWR.n296 VPWR.n266 0.120292
R439 VPWR.n296 VPWR.n295 0.120292
R440 VPWR.n295 VPWR.n294 0.120292
R441 VPWR.n294 VPWR.n268 0.120292
R442 VPWR.n289 VPWR.n268 0.120292
R443 VPWR.n289 VPWR.n288 0.120292
R444 VPWR.n288 VPWR.n287 0.120292
R445 VPWR.n287 VPWR.n271 0.120292
R446 VPWR.n283 VPWR.n271 0.120292
R447 VPWR.n283 VPWR.n282 0.120292
R448 VPWR.n282 VPWR.n274 0.120292
R449 VPWR.n278 VPWR.n274 0.120292
R450 VPWR.n220 VPWR.n219 0.12023
R451 VPWR.n166 VPWR.n165 0.12023
R452 VPWR.n219 VPWR.n218 0.119565
R453 VPWR.n167 VPWR.n166 0.119565
R454 VPWR.n228 VPWR.n227 0.118556
R455 VPWR.n147 VPWR.n87 0.118474
R456 VPWR.n104 VPWR.n103 0.117381
R457 VPWR.n197 VPWR.n196 0.117018
R458 VPWR.n198 VPWR.n197 0.116571
R459 VPWR.n218 VPWR.n217 0.115278
R460 VPWR.n168 VPWR.n167 0.115278
R461 VPWR.n227 VPWR.n11 0.114758
R462 VPWR.n90 VPWR.n89 0.114696
R463 VPWR.n207 VPWR.n29 0.114511
R464 VPWR.n217 VPWR.n216 0.114352
R465 VPWR.n169 VPWR.n168 0.114352
R466 VPWR.n102 VPWR.n101 0.114094
R467 VPWR.n216 VPWR.n215 0.113756
R468 VPWR.n170 VPWR.n169 0.113235
R469 VPWR.n92 VPWR.n91 0.113192
R470 VPWR.n101 VPWR.n100 0.113154
R471 VPWR.n91 VPWR.n90 0.112678
R472 VPWR.n94 VPWR.n93 0.112433
R473 VPWR.n209 VPWR.n208 0.112207
R474 VPWR.n199 VPWR.n198 0.111422
R475 VPWR.n215 VPWR.n214 0.111333
R476 VPWR.n98 VPWR.n97 0.111285
R477 VPWR.n214 VPWR.n213 0.111081
R478 VPWR.n172 VPWR.n171 0.111081
R479 VPWR.n12 VPWR.n11 0.111077
R480 VPWR.n171 VPWR.n170 0.110429
R481 VPWR.n96 VPWR.n95 0.110229
R482 VPWR.n173 VPWR.n172 0.11011
R483 VPWR.n93 VPWR.n92 0.109923
R484 VPWR.n103 VPWR.n102 0.10979
R485 VPWR.n201 VPWR.n200 0.109555
R486 VPWR.n183 VPWR.n182 0.108951
R487 VPWR.n211 VPWR.n210 0.108673
R488 VPWR.n175 VPWR.n174 0.108673
R489 VPWR.n213 VPWR.n212 0.108622
R490 VPWR.n99 VPWR.n98 0.108359
R491 VPWR.n100 VPWR.n99 0.108286
R492 VPWR.n95 VPWR.n94 0.10823
R493 VPWR.n200 VPWR.n199 0.107819
R494 VPWR.n97 VPWR.n96 0.107643
R495 VPWR.n236 VPWR.n235 0.107643
R496 VPWR.n212 VPWR.n211 0.107267
R497 VPWR.n174 VPWR.n173 0.107267
R498 VPWR.n177 VPWR.n176 0.107106
R499 VPWR.n13 VPWR.n12 0.106561
R500 VPWR.n202 VPWR.n201 0.105203
R501 VPWR.n203 VPWR.n202 0.105131
R502 VPWR.n182 VPWR.n181 0.104693
R503 VPWR.n205 VPWR.n204 0.104583
R504 VPWR.n181 VPWR.n180 0.104583
R505 VPWR.n204 VPWR.n203 0.104127
R506 VPWR.n206 VPWR.n205 0.103965
R507 VPWR.n180 VPWR.n179 0.103965
R508 VPWR.n207 VPWR.n206 0.103813
R509 VPWR.n179 VPWR.n178 0.103813
R510 VPWR.n178 VPWR.n177 0.103788
R511 VPWR.n210 VPWR.n209 0.103439
R512 VPWR.n176 VPWR.n175 0.103439
R513 VPWR.n223 VPWR.n222 0.100519
R514 VPWR VPWR.n0 0.0981562
R515 VPWR VPWR.n337 0.0981562
R516 VPWR.n302 VPWR 0.0981562
R517 VPWR.n15 VPWR.n14 0.0979265
R518 VPWR.n79 VPWR.n78 0.0979265
R519 VPWR.n16 VPWR.n15 0.0960882
R520 VPWR.n78 VPWR.n77 0.0960882
R521 VPWR.n17 VPWR.n16 0.0915714
R522 VPWR.n77 VPWR.n76 0.0915714
R523 VPWR.n18 VPWR.n17 0.088
R524 VPWR.n76 VPWR.n75 0.088
R525 VPWR.n19 VPWR.n18 0.0855694
R526 VPWR.n75 VPWR.n74 0.0855694
R527 VPWR.n146 VPWR.n88 0.0849982
R528 VPWR.n223 VPWR.n13 0.0844552
R529 VPWR.n230 VPWR.n229 0.0832089
R530 VPWR VPWR.n341 0.0825312
R531 VPWR VPWR.n307 0.0825312
R532 VPWR.n20 VPWR.n19 0.0820972
R533 VPWR.n74 VPWR.n73 0.0820972
R534 VPWR.n21 VPWR.n20 0.0792671
R535 VPWR.n73 VPWR.n72 0.0792671
R536 VPWR.n22 VPWR.n21 0.0775548
R537 VPWR.n72 VPWR.n71 0.0765135
R538 VPWR.n146 VPWR.n145 0.0741301
R539 VPWR.n71 VPWR.n70 0.0731351
R540 VPWR.n145 VPWR.n144 0.0724178
R541 VPWR.n23 VPWR.n22 0.0721667
R542 VPWR.n24 VPWR.n23 0.0705
R543 VPWR.n70 VPWR.n69 0.0705
R544 VPWR.n144 VPWR.n143 0.0688333
R545 VPWR.n25 VPWR.n24 0.0679342
R546 VPWR.n69 VPWR.n68 0.0679342
R547 VPWR.n29 VPWR.n28 0.0676642
R548 VPWR.n143 VPWR.n142 0.0655
R549 VPWR.n26 VPWR.n25 0.0646447
R550 VPWR.n68 VPWR.n67 0.0646447
R551 VPWR.n142 VPWR.n141 0.0646447
R552 VPWR.n27 VPWR.n26 0.063
R553 VPWR.n67 VPWR.n66 0.063
R554 VPWR.n343 VPWR 0.0603958
R555 VPWR VPWR.n342 0.0603958
R556 VPWR.n341 VPWR 0.0603958
R557 VPWR.n338 VPWR 0.0603958
R558 VPWR.n311 VPWR 0.0603958
R559 VPWR.n308 VPWR 0.0603958
R560 VPWR.n307 VPWR 0.0603958
R561 VPWR VPWR.n306 0.0603958
R562 VPWR.n141 VPWR.n140 0.0597105
R563 VPWR.n28 VPWR.n27 0.0589416
R564 VPWR.n66 VPWR.n65 0.0589416
R565 VPWR.n140 VPWR.n139 0.0581923
R566 VPWR.n65 VPWR.n64 0.057462
R567 VPWR.n154 VPWR 0.0573182
R568 VPWR.n83 VPWR 0.0573182
R569 VPWR.n81 VPWR 0.0573182
R570 VPWR.n54 VPWR 0.0573182
R571 VPWR.n31 VPWR 0.0573182
R572 VPWR.n10 VPWR 0.0573182
R573 VPWR.n7 VPWR 0.0573182
R574 VPWR.n4 VPWR 0.0573182
R575 VPWR.n57 VPWR 0.0573182
R576 VPWR.n160 VPWR 0.0573182
R577 VPWR.n139 VPWR.n138 0.0556948
R578 VPWR.n64 VPWR.n63 0.0542975
R579 VPWR.n33 VPWR.n32 0.0527152
R580 VPWR.n63 VPWR.n62 0.0527152
R581 VPWR.n138 VPWR.n137 0.0527152
R582 VPWR.n115 VPWR 0.0505
R583 VPWR.n149 VPWR 0.0505
R584 VPWR.n86 VPWR 0.0505
R585 VPWR.n110 VPWR 0.0505
R586 VPWR.n123 VPWR 0.0505
R587 VPWR.n120 VPWR 0.0505
R588 VPWR.n137 VPWR.n136 0.0495506
R589 VPWR.n34 VPWR.n33 0.0483395
R590 VPWR.n62 VPWR.n61 0.0483395
R591 VPWR.n136 VPWR.n135 0.0479684
R592 VPWR.n35 VPWR.n34 0.047375
R593 VPWR.n61 VPWR.n60 0.047375
R594 VPWR.n32 VPWR.n29 0.0472033
R595 VPWR.n60 VPWR.n59 0.0463861
R596 VPWR.n36 VPWR.n35 0.0452531
R597 VPWR.n135 VPWR.n134 0.0452531
R598 VPWR.n134 VPWR.n133 0.0426875
R599 VPWR.n37 VPWR.n36 0.0416585
R600 VPWR.n59 VPWR.n58 0.0406786
R601 VPWR.n88 VPWR.n87 0.039507
R602 VPWR.n133 VPWR.n132 0.0390802
R603 VPWR.n38 VPWR.n37 0.0386098
R604 VPWR.n39 VPWR.n38 0.0386098
R605 VPWR.n132 VPWR.n131 0.0386098
R606 VPWR.n342 VPWR 0.0382604
R607 VPWR.n308 VPWR 0.0382604
R608 VPWR.n131 VPWR.n130 0.035561
R609 VPWR.n40 VPWR.n39 0.0351386
R610 VPWR.n126 VPWR.n125 0.0350681
R611 VPWR.n130 VPWR.n129 0.0325122
R612 VPWR.n41 VPWR.n40 0.0321265
R613 VPWR.n129 VPWR.n128 0.0306205
R614 VPWR.n42 VPWR.n41 0.0302619
R615 VPWR.n128 VPWR.n127 0.0276084
R616 VPWR.n43 VPWR.n42 0.0272857
R617 VPWR.n44 VPWR.n43 0.0257976
R618 VPWR.n127 VPWR.n126 0.0257976
R619 VPWR.n55 VPWR.n52 0.0244583
R620 VPWR.n45 VPWR.n44 0.0243095
R621 VPWR.n236 VPWR.n1 0.0243095
R622 VPWR.n185 VPWR.n55 0.0239375
R623 VPWR.n184 VPWR.n58 0.0227865
R624 VPWR.n338 VPWR 0.0226354
R625 VPWR.n306 VPWR 0.0226354
R626 VPWR VPWR.n373 0.0224072
R627 VPWR.n2 VPWR.n1 0.0214028
R628 VPWR.n46 VPWR.n45 0.0210882
R629 VPWR.n47 VPWR.n46 0.0198452
R630 VPWR.n48 VPWR.n47 0.0166765
R631 VPWR.n49 VPWR.n48 0.0152059
R632 VPWR.n234 VPWR.n233 0.01479
R633 VPWR.n111 VPWR.n108 0.0131488
R634 VPWR.n234 VPWR.n1 0.0124293
R635 VPWR.n50 VPWR.n49 0.0121279
R636 VPWR.n51 VPWR.n50 0.0107941
R637 VPWR.n162 VPWR.n161 0.0104434
R638 VPWR.n52 VPWR.n51 0.00785294
R639 VPWR.n229 VPWR.n228 0.00590163
R640 VGND.n439 VGND.n62 171881
R641 VGND.n457 VGND.n456 156689
R642 VGND.n65 VGND.t67 151322
R643 VGND.n436 VGND.n229 130569
R644 VGND.n483 VGND.n482 130542
R645 VGND.n272 VGND.n226 49690.4
R646 VGND.n280 VGND.n3 48636.9
R647 VGND.n442 VGND.n229 45450.3
R648 VGND.n484 VGND.n483 44132.5
R649 VGND.n436 VGND.n435 44106
R650 VGND.n437 VGND.n231 43377.2
R651 VGND.n435 VGND.t16 31560.8
R652 VGND.n485 VGND.n484 30151.8
R653 VGND.n435 VGND.n231 29891.4
R654 VGND.n484 VGND.n1 29891.4
R655 VGND.n304 VGND.t65 18687.3
R656 VGND.n442 VGND.n62 16600.2
R657 VGND.n290 VGND.n285 16072.7
R658 VGND.n230 VGND.n61 14081.5
R659 VGND.n307 VGND.n272 13406.4
R660 VGND.n304 VGND.n303 13301.5
R661 VGND.n275 VGND.n274 12272.6
R662 VGND.n298 VGND.n275 12077.4
R663 VGND.n443 VGND.n442 11373.6
R664 VGND.n437 VGND.n436 10649.3
R665 VGND.n483 VGND.n3 10649.2
R666 VGND.n442 VGND.n226 8289.38
R667 VGND.n277 VGND.n275 6135.59
R668 VGND.n438 VGND.n437 6127.89
R669 VGND.n304 VGND 5326.64
R670 VGND.n307 VGND.n273 4245.54
R671 VGND.t12 VGND.n289 4169.04
R672 VGND.n434 VGND.n228 4044.64
R673 VGND.t37 VGND.n228 3942.35
R674 VGND.n442 VGND.n227 3472.59
R675 VGND.n456 VGND.n455 3462.51
R676 VGND.n289 VGND.n288 3164.24
R677 VGND.n291 VGND.n290 3164.24
R678 VGND.n290 VGND.n287 3154.4
R679 VGND.n277 VGND.n276 3108.35
R680 VGND.n280 VGND.n277 3022.83
R681 VGND.n289 VGND.n285 2949.38
R682 VGND.n274 VGND.n230 2758.39
R683 VGND.n442 VGND.n441 2554.5
R684 VGND.n455 VGND.t29 2387.95
R685 VGND.n304 VGND 2380.9
R686 VGND.n299 VGND.n230 2252.33
R687 VGND.n442 VGND.n438 2096.68
R688 VGND.n307 VGND.n306 1953.47
R689 VGND.n457 VGND.n62 1821.62
R690 VGND.n279 VGND.t80 1524.56
R691 VGND.n313 VGND.n231 1397.72
R692 VGND.n303 VGND.t6 1303.08
R693 VGND.n281 VGND.n280 1261.32
R694 VGND.n434 VGND.n433 1170
R695 VGND.n303 VGND.n302 1170
R696 VGND.n449 VGND.n64 1170
R697 VGND.n220 VGND.n63 1170
R698 VGND.n454 VGND.n453 1170
R699 VGND.n441 VGND.n440 1170
R700 VGND.n459 VGND.n458 1170
R701 VGND.n445 VGND.n444 1170
R702 VGND.n377 VGND.n227 1170
R703 VGND.n306 VGND.n305 1170
R704 VGND.n309 VGND.n308 1170
R705 VGND.n297 VGND.n296 1170
R706 VGND.n287 VGND.n286 1170
R707 VGND.n279 VGND.n278 1170
R708 VGND.n481 VGND.n480 1170
R709 VGND.n24 VGND.n2 1170
R710 VGND.n282 VGND.n281 1170
R711 VGND.n487 VGND.n486 1170
R712 VGND.n481 VGND.t14 1134.17
R713 VGND.n307 VGND.n299 1052.01
R714 VGND.t23 VGND.n457 876.702
R715 VGND.n229 VGND.t41 844.357
R716 VGND.n61 VGND.n4 843.24
R717 VGND.t32 VGND.n485 753.322
R718 VGND.n273 VGND.n231 747.253
R719 VGND.t67 VGND.n63 713.466
R720 VGND.t71 VGND.n1 696.106
R721 VGND.n455 VGND.n64 634.212
R722 VGND.t2 VGND.n231 629.832
R723 VGND.n300 VGND 589.678
R724 VGND.n300 VGND 589.678
R725 VGND.n485 VGND.n2 585.742
R726 VGND.n486 VGND.n1 546.058
R727 VGND.t29 VGND.n454 508.485
R728 VGND.n442 VGND.n228 493.118
R729 VGND.n273 VGND.t48 467.337
R730 VGND.t16 VGND.n434 380.034
R731 VGND.n444 VGND.n443 333.548
R732 VGND.n285 VGND.t51 302.156
R733 VGND.n487 VGND.t33 282.339
R734 VGND.n24 VGND.t15 282.339
R735 VGND.n480 VGND.t28 282.339
R736 VGND.n459 VGND.t24 282.339
R737 VGND.n440 VGND.t26 282.339
R738 VGND.n286 VGND.t70 282.339
R739 VGND.n296 VGND.t76 282.339
R740 VGND.n278 VGND.t81 282.339
R741 VGND.n282 VGND.t72 282.339
R742 VGND.n288 VGND.t74 282.339
R743 VGND.n453 VGND.t30 282.339
R744 VGND.n433 VGND.t17 282.339
R745 VGND.n305 VGND.t3 282.339
R746 VGND.n309 VGND.t52 282.339
R747 VGND.n291 VGND.t13 282.339
R748 VGND.n313 VGND.t49 282.339
R749 VGND.n302 VGND.t7 282.339
R750 VGND.n377 VGND.t42 282.339
R751 VGND.n445 VGND.t45 282.339
R752 VGND.n449 VGND.t5 282.339
R753 VGND.n220 VGND.t68 282.339
R754 VGND.t41 VGND.n227 266.457
R755 VGND.n119 VGND.t56 251
R756 VGND.n153 VGND.t78 251
R757 VGND.n187 VGND.t40 251
R758 VGND.t25 VGND.n439 248.936
R759 VGND.n106 VGND.t11 243.028
R760 VGND.n140 VGND.t62 243.028
R761 VGND.n174 VGND.t22 243.028
R762 VGND.n289 VGND.t73 236.923
R763 VGND.n307 VGND.n304 219.505
R764 VGND.n93 VGND.n92 218.506
R765 VGND.n80 VGND.n79 218.506
R766 VGND.n189 VGND.n188 218.506
R767 VGND.n280 VGND.n279 212.281
R768 VGND.n297 VGND.n276 204.773
R769 VGND.n90 VGND.n89 200.201
R770 VGND.n77 VGND.n76 200.201
R771 VGND.n197 VGND.n196 200.201
R772 VGND.n102 VGND.n101 199.739
R773 VGND.n136 VGND.n135 199.739
R774 VGND.n170 VGND.n169 199.739
R775 VGND.n112 VGND.n98 199.53
R776 VGND.n146 VGND.n85 199.53
R777 VGND.n180 VGND.n72 199.53
R778 VGND.n454 VGND.n65 190.542
R779 VGND.n441 VGND.t25 187.446
R780 VGND.n298 VGND.t75 183.096
R781 VGND.n486 VGND.t32 170.459
R782 VGND.n306 VGND.t2 169.868
R783 VGND.t14 VGND.n2 166.094
R784 VGND.n304 VGND.n228 165.339
R785 VGND.n442 VGND.t44 159.488
R786 VGND.n281 VGND.t71 158.115
R787 VGND.n456 VGND.n63 144.5
R788 VGND.t75 VGND.n297 140.434
R789 VGND.n443 VGND.t4 132.02
R790 VGND.t0 VGND.n226 128.904
R791 VGND.n458 VGND.t23 124.144
R792 VGND.n444 VGND.t44 122.326
R793 VGND.t69 VGND.n285 120.314
R794 VGND.n308 VGND.t51 111.326
R795 VGND.n299 VGND.n298 104.849
R796 VGND VGND.t43 102.412
R797 VGND.t4 VGND.n64 101.258
R798 VGND.n482 VGND.n4 100.996
R799 VGND.t10 VGND.n272 94.8614
R800 VGND.t55 VGND.t19 93.0774
R801 VGND.n287 VGND.t69 92.2804
R802 VGND.n98 VGND.t20 74.8666
R803 VGND.n85 VGND.t36 74.8666
R804 VGND.n72 VGND.t47 74.8666
R805 VGND.n290 VGND.t12 55.9751
R806 VGND.n89 VGND.t59 54.2862
R807 VGND.n76 VGND.t77 54.2862
R808 VGND.n196 VGND.t38 54.2862
R809 VGND.n482 VGND.n481 46.6396
R810 VGND VGND.t66 45.7764
R811 VGND.n274 VGND.n3 45.2738
R812 VGND.n458 VGND.n61 40.8576
R813 VGND.n98 VGND.t63 40.0005
R814 VGND.n85 VGND.t82 40.0005
R815 VGND.n72 VGND.t34 40.0005
R816 VGND.n101 VGND.t21 38.5719
R817 VGND.n101 VGND.t64 38.5719
R818 VGND.n135 VGND.t9 38.5719
R819 VGND.n135 VGND.t61 38.5719
R820 VGND.n169 VGND.t54 38.5719
R821 VGND.n169 VGND.t53 38.5719
R822 VGND.n308 VGND.n307 36.639
R823 VGND.n108 VGND.n107 34.6358
R824 VGND.n108 VGND.n97 34.6358
R825 VGND.n114 VGND.n113 34.6358
R826 VGND.n114 VGND.n95 34.6358
R827 VGND.n118 VGND.n95 34.6358
R828 VGND.n124 VGND.n123 34.6358
R829 VGND.n125 VGND.n124 34.6358
R830 VGND.n130 VGND.n129 34.6358
R831 VGND.n130 VGND.n88 34.6358
R832 VGND.n134 VGND.n88 34.6358
R833 VGND.n142 VGND.n141 34.6358
R834 VGND.n142 VGND.n84 34.6358
R835 VGND.n148 VGND.n147 34.6358
R836 VGND.n148 VGND.n82 34.6358
R837 VGND.n152 VGND.n82 34.6358
R838 VGND.n158 VGND.n157 34.6358
R839 VGND.n159 VGND.n158 34.6358
R840 VGND.n164 VGND.n163 34.6358
R841 VGND.n164 VGND.n75 34.6358
R842 VGND.n168 VGND.n75 34.6358
R843 VGND.n176 VGND.n175 34.6358
R844 VGND.n176 VGND.n71 34.6358
R845 VGND.n182 VGND.n181 34.6358
R846 VGND.n182 VGND.n69 34.6358
R847 VGND.n186 VGND.n69 34.6358
R848 VGND.n194 VGND.n67 34.6358
R849 VGND.n195 VGND.n194 34.6358
R850 VGND.n120 VGND.n93 32.7534
R851 VGND.n154 VGND.n80 32.7534
R852 VGND.n190 VGND.n189 32.7534
R853 VGND.n120 VGND.n119 31.2476
R854 VGND.n154 VGND.n153 31.2476
R855 VGND.n190 VGND.n187 31.2476
R856 VGND.n112 VGND.n97 30.8711
R857 VGND.n146 VGND.n84 30.8711
R858 VGND.n180 VGND.n71 30.8711
R859 VGND.n107 VGND.n106 27.4829
R860 VGND.n141 VGND.n140 27.4829
R861 VGND.n175 VGND.n174 27.4829
R862 VGND.t8 VGND.t35 27.1458
R863 VGND.n89 VGND.t50 25.9346
R864 VGND.n76 VGND.t46 25.9346
R865 VGND.n196 VGND.t18 25.9346
R866 VGND.t65 VGND.t55 25.3851
R867 VGND.n92 VGND.t60 24.9236
R868 VGND.n92 VGND.t58 24.9236
R869 VGND.n79 VGND.t1 24.9236
R870 VGND.n79 VGND.t79 24.9236
R871 VGND.n188 VGND.t31 24.9236
R872 VGND.n188 VGND.t39 24.9236
R873 VGND.n125 VGND.n90 23.7181
R874 VGND.n159 VGND.n77 23.7181
R875 VGND.n197 VGND.n195 23.7181
R876 VGND.n102 VGND.n100 22.9652
R877 VGND.n106 VGND.n100 22.9652
R878 VGND.n136 VGND.n87 22.9652
R879 VGND.n140 VGND.n87 22.9652
R880 VGND.n170 VGND.n74 22.9652
R881 VGND.n174 VGND.n74 22.9652
R882 VGND.n119 VGND.n118 22.2123
R883 VGND.n153 VGND.n152 22.2123
R884 VGND.n187 VGND.n186 22.2123
R885 VGND.n129 VGND.n90 21.4593
R886 VGND.n136 VGND.n134 21.4593
R887 VGND.n163 VGND.n77 21.4593
R888 VGND.n170 VGND.n168 21.4593
R889 VGND.n295 VGND.n284 20.9265
R890 VGND.n285 VGND.n276 20.0607
R891 VGND.t0 VGND.t37 19.8983
R892 VGND.t0 VGND.n300 19.7425
R893 VGND.n218 VGND 17.3883
R894 VGND.n461 VGND.n60 17.0502
R895 VGND.n438 VGND.n230 14.7835
R896 VGND.n433 VGND.n432 13.3141
R897 VGND.n305 VGND.n252 13.3141
R898 VGND.n310 VGND.n309 13.3141
R899 VGND.n292 VGND.n291 13.3141
R900 VGND.n314 VGND.n313 13.3141
R901 VGND.n302 VGND.n301 13.3141
R902 VGND.n378 VGND.n377 13.3141
R903 VGND.n446 VGND.n445 13.3141
R904 VGND.n450 VGND.n449 13.3141
R905 VGND.n221 VGND.n220 13.3141
R906 VGND VGND.n24 13.2586
R907 VGND.n480 VGND 13.2586
R908 VGND VGND.n459 13.2586
R909 VGND.n440 VGND 13.2586
R910 VGND.n286 VGND 13.2586
R911 VGND.n296 VGND 13.2586
R912 VGND.n278 VGND 13.2586
R913 VGND VGND.n282 13.2586
R914 VGND.n288 VGND 13.2586
R915 VGND.n453 VGND 13.2586
R916 VGND VGND.n487 13.2586
R917 VGND VGND.n60 10.8878
R918 VGND.n113 VGND.n112 10.5417
R919 VGND.n147 VGND.n146 10.5417
R920 VGND.n181 VGND.n180 10.5417
R921 VGND.n451 VGND.n448 9.52816
R922 VGND VGND.n452 9.46719
R923 VGND.n104 VGND.n100 9.3005
R924 VGND.n106 VGND.n105 9.3005
R925 VGND.n107 VGND.n99 9.3005
R926 VGND.n109 VGND.n108 9.3005
R927 VGND.n110 VGND.n97 9.3005
R928 VGND.n112 VGND.n111 9.3005
R929 VGND.n113 VGND.n96 9.3005
R930 VGND.n115 VGND.n114 9.3005
R931 VGND.n116 VGND.n95 9.3005
R932 VGND.n118 VGND.n117 9.3005
R933 VGND.n119 VGND.n94 9.3005
R934 VGND.n121 VGND.n120 9.3005
R935 VGND.n123 VGND.n122 9.3005
R936 VGND.n124 VGND.n91 9.3005
R937 VGND.n126 VGND.n125 9.3005
R938 VGND.n127 VGND.n90 9.3005
R939 VGND.n129 VGND.n128 9.3005
R940 VGND.n131 VGND.n130 9.3005
R941 VGND.n132 VGND.n88 9.3005
R942 VGND.n134 VGND.n133 9.3005
R943 VGND.n137 VGND.n136 9.3005
R944 VGND.n138 VGND.n87 9.3005
R945 VGND.n140 VGND.n139 9.3005
R946 VGND.n141 VGND.n86 9.3005
R947 VGND.n143 VGND.n142 9.3005
R948 VGND.n144 VGND.n84 9.3005
R949 VGND.n146 VGND.n145 9.3005
R950 VGND.n147 VGND.n83 9.3005
R951 VGND.n149 VGND.n148 9.3005
R952 VGND.n150 VGND.n82 9.3005
R953 VGND.n152 VGND.n151 9.3005
R954 VGND.n153 VGND.n81 9.3005
R955 VGND.n155 VGND.n154 9.3005
R956 VGND.n157 VGND.n156 9.3005
R957 VGND.n158 VGND.n78 9.3005
R958 VGND.n160 VGND.n159 9.3005
R959 VGND.n161 VGND.n77 9.3005
R960 VGND.n163 VGND.n162 9.3005
R961 VGND.n165 VGND.n164 9.3005
R962 VGND.n166 VGND.n75 9.3005
R963 VGND.n168 VGND.n167 9.3005
R964 VGND.n171 VGND.n170 9.3005
R965 VGND.n172 VGND.n74 9.3005
R966 VGND.n174 VGND.n173 9.3005
R967 VGND.n175 VGND.n73 9.3005
R968 VGND.n177 VGND.n176 9.3005
R969 VGND.n178 VGND.n71 9.3005
R970 VGND.n180 VGND.n179 9.3005
R971 VGND.n181 VGND.n70 9.3005
R972 VGND.n183 VGND.n182 9.3005
R973 VGND.n184 VGND.n69 9.3005
R974 VGND.n186 VGND.n185 9.3005
R975 VGND.n187 VGND.n68 9.3005
R976 VGND.n191 VGND.n190 9.3005
R977 VGND.n192 VGND.n67 9.3005
R978 VGND.n194 VGND.n193 9.3005
R979 VGND.n195 VGND.n66 9.3005
R980 VGND.n293 VGND.n292 9.16992
R981 VGND VGND.n295 8.69654
R982 VGND.n311 VGND.n310 8.60727
R983 VGND.n460 VGND 8.50779
R984 VGND.n312 VGND.n311 8.47796
R985 VGND.n222 VGND.n221 7.73586
R986 VGND.n294 VGND 7.66873
R987 VGND.t43 VGND.t8 7.40375
R988 VGND VGND.n479 7.24133
R989 VGND.n315 VGND.n314 7.18609
R990 VGND.n103 VGND.n102 7.12576
R991 VGND.n198 VGND.n197 7.12063
R992 VGND.n451 VGND.n450 6.8256
R993 VGND VGND.n271 6.67637
R994 VGND.n447 VGND.n446 6.61112
R995 VGND.n334 VGND.n252 6.60276
R996 VGND.n25 VGND 6.5915
R997 VGND VGND.n0 6.55995
R998 VGND.n284 VGND 6.30778
R999 VGND.n411 VGND.n378 6.21471
R1000 VGND.n283 VGND 6.20286
R1001 VGND.n301 VGND.n232 6.13644
R1002 VGND.n432 VGND.n431 5.99894
R1003 VGND.t19 VGND.t57 4.23127
R1004 VGND.n311 VGND.n271 3.52873
R1005 VGND.n219 VGND 3.40017
R1006 VGND.t66 VGND.t10 3.3096
R1007 VGND.n219 VGND.n218 3.28674
R1008 VGND.n284 VGND.n283 2.92676
R1009 VGND.n452 VGND.n451 2.38171
R1010 VGND.n439 VGND.n65 2.10058
R1011 VGND.n4 VGND.t27 1.91332
R1012 VGND.n123 VGND.n93 1.88285
R1013 VGND.n157 VGND.n80 1.88285
R1014 VGND.n189 VGND.n67 1.88285
R1015 VGND.n295 VGND.n294 1.59945
R1016 VGND.n283 VGND.n0 1.28972
R1017 VGND.t35 VGND.t0 1.23438
R1018 VGND.n223 VGND.n219 1.1273
R1019 VGND.n294 VGND.n293 1.05629
R1020 VGND.n452 VGND.n223 0.953601
R1021 VGND.n293 VGND.n271 0.951859
R1022 VGND.n199 uo_out[4] 0.844933
R1023 VGND.n222 VGND.n60 0.753637
R1024 VGND.n26 VGND.n0 0.663554
R1025 VGND.n218 VGND.n217 0.646593
R1026 VGND.n202 VGND.n201 0.5786
R1027 VGND.n200 VGND.n199 0.577033
R1028 VGND.n201 VGND.n200 0.577033
R1029 VGND.n204 VGND.n203 0.577033
R1030 VGND.n205 VGND.n204 0.577033
R1031 VGND.n206 VGND.n205 0.577033
R1032 VGND.n207 VGND.n206 0.577033
R1033 VGND.n208 VGND.n207 0.577033
R1034 VGND.n209 VGND.n208 0.577033
R1035 VGND.n210 VGND.n209 0.577033
R1036 VGND.n211 VGND.n210 0.577033
R1037 VGND.n212 VGND.n211 0.577033
R1038 VGND.n213 VGND.n212 0.577033
R1039 VGND.n214 VGND.n213 0.577033
R1040 VGND.n215 VGND.n214 0.577033
R1041 VGND.n216 VGND.n215 0.577033
R1042 VGND.n217 VGND.n216 0.577033
R1043 VGND.n203 VGND.n202 0.575467
R1044 VGND.n357 VGND.n356 0.457033
R1045 VGND.n354 VGND.n232 0.297375
R1046 VGND.n217 uio_oe[7] 0.2684
R1047 VGND.n199 uo_out[5] 0.2684
R1048 VGND.n200 uo_out[6] 0.2684
R1049 VGND.n201 uo_out[7] 0.2684
R1050 VGND.n202 uio_out[0] 0.2684
R1051 VGND.n203 uio_out[1] 0.2684
R1052 VGND.n204 uio_out[2] 0.2684
R1053 VGND.n205 uio_out[3] 0.2684
R1054 VGND.n206 uio_out[4] 0.2684
R1055 VGND.n207 uio_out[5] 0.2684
R1056 VGND.n208 uio_out[6] 0.2684
R1057 VGND.n209 uio_out[7] 0.2684
R1058 VGND.n210 uio_oe[0] 0.2684
R1059 VGND.n211 uio_oe[1] 0.2684
R1060 VGND.n212 uio_oe[2] 0.2684
R1061 VGND.n213 uio_oe[3] 0.2684
R1062 VGND.n214 uio_oe[4] 0.2684
R1063 VGND.n215 uio_oe[5] 0.2684
R1064 VGND.n216 uio_oe[6] 0.2684
R1065 VGND.n354 VGND.n353 0.240747
R1066 VGND.n43 VGND.n7 0.232444
R1067 VGND.n353 VGND.n352 0.201889
R1068 VGND.n352 VGND.n351 0.183192
R1069 VGND.n448 VGND.n224 0.181207
R1070 VGND.n27 VGND.n26 0.177735
R1071 VGND.n315 VGND.n312 0.15732
R1072 VGND.n462 VGND.n461 0.155253
R1073 VGND VGND.n198 0.152603
R1074 VGND.n44 VGND.n43 0.152388
R1075 VGND.n198 VGND.n66 0.148519
R1076 VGND.n350 VGND.n349 0.145639
R1077 VGND.n411 VGND.n410 0.14536
R1078 VGND.n351 VGND.n350 0.14425
R1079 VGND.n104 VGND.n103 0.143396
R1080 VGND.n353 VGND.n233 0.135917
R1081 VGND.n355 VGND.n354 0.135115
R1082 VGND.n351 VGND.n235 0.134528
R1083 VGND.n352 VGND.n234 0.133742
R1084 VGND.n356 VGND.n232 0.133539
R1085 VGND.n349 VGND.n237 0.133139
R1086 VGND.n350 VGND.n236 0.133139
R1087 VGND.n348 VGND.n238 0.13175
R1088 VGND.n28 VGND.n22 0.131182
R1089 VGND.n345 VGND.n241 0.131118
R1090 VGND.n347 VGND.n239 0.131056
R1091 VGND.n346 VGND.n240 0.130361
R1092 VGND.n341 VGND.n245 0.129761
R1093 VGND.n30 VGND.n20 0.129761
R1094 VGND.n344 VGND.n242 0.129713
R1095 VGND.n27 VGND.n23 0.129713
R1096 VGND.n31 VGND.n19 0.128341
R1097 VGND.n342 VGND.n244 0.128309
R1098 VGND.n29 VGND.n21 0.128309
R1099 VGND.n343 VGND.n243 0.128278
R1100 VGND.n36 VGND.n14 0.12768
R1101 VGND.n34 VGND.n16 0.127655
R1102 VGND.n339 VGND.n247 0.127631
R1103 VGND.n430 VGND.n358 0.127631
R1104 VGND.n32 VGND.n18 0.127631
R1105 VGND.n37 VGND.n13 0.126953
R1106 VGND.n35 VGND.n15 0.126937
R1107 VGND.n338 VGND.n248 0.12692
R1108 VGND.n429 VGND.n359 0.12692
R1109 VGND.n33 VGND.n17 0.12692
R1110 VGND.n340 VGND.n246 0.126904
R1111 VGND.n397 VGND.n392 0.126368
R1112 VGND.n462 VGND.n59 0.126345
R1113 VGND.n464 VGND.n57 0.126333
R1114 VGND.n466 VGND.n55 0.126322
R1115 VGND.n468 VGND.n53 0.126312
R1116 VGND.n42 VGND.n8 0.126244
R1117 VGND.n335 VGND.n251 0.126218
R1118 VGND.n426 VGND.n362 0.126218
R1119 VGND.n337 VGND.n249 0.12621
R1120 VGND.n428 VGND.n360 0.12621
R1121 VGND.n331 VGND.n255 0.1255
R1122 VGND.n332 VGND.n254 0.1255
R1123 VGND.n333 VGND.n253 0.1255
R1124 VGND.n336 VGND.n250 0.1255
R1125 VGND.n427 VGND.n361 0.1255
R1126 VGND.n425 VGND.n363 0.1255
R1127 VGND.n424 VGND.n364 0.1255
R1128 VGND.n423 VGND.n365 0.1255
R1129 VGND.n38 VGND.n12 0.1255
R1130 VGND.n39 VGND.n11 0.1255
R1131 VGND.n40 VGND.n10 0.1255
R1132 VGND.n473 VGND.n48 0.1255
R1133 VGND.n471 VGND.n50 0.1255
R1134 VGND.n463 VGND.n58 0.1255
R1135 VGND.n328 VGND.n258 0.124765
R1136 VGND.n420 VGND.n368 0.124765
R1137 VGND.n41 VGND.n9 0.124765
R1138 VGND.n479 VGND.n478 0.124747
R1139 VGND.n476 VGND.n45 0.124738
R1140 VGND.n474 VGND.n47 0.124728
R1141 VGND.n470 VGND.n51 0.124709
R1142 VGND.n405 VGND.n384 0.124688
R1143 VGND.n403 VGND.n386 0.124678
R1144 VGND.n401 VGND.n388 0.124667
R1145 VGND.n399 VGND.n390 0.124655
R1146 VGND.n398 VGND.n391 0.124655
R1147 VGND.n396 VGND.n393 0.124644
R1148 VGND.n330 VGND.n256 0.124047
R1149 VGND.n422 VGND.n366 0.124047
R1150 VGND.n326 VGND.n260 0.124012
R1151 VGND.n418 VGND.n370 0.124012
R1152 VGND.n324 VGND.n262 0.123994
R1153 VGND.n416 VGND.n372 0.123994
R1154 VGND.n477 VGND.n6 0.123994
R1155 VGND.n475 VGND.n46 0.123976
R1156 VGND.n318 VGND.n268 0.123938
R1157 VGND.n316 VGND.n270 0.123918
R1158 VGND.n408 VGND.n381 0.123918
R1159 VGND.n469 VGND.n52 0.123918
R1160 VGND.n467 VGND.n54 0.123897
R1161 VGND.n465 VGND.n56 0.123877
R1162 VGND.n400 VGND.n389 0.123833
R1163 VGND.n410 VGND.n409 0.123779
R1164 VGND.n329 VGND.n257 0.12332
R1165 VGND.n421 VGND.n367 0.12332
R1166 VGND.n327 VGND.n259 0.123294
R1167 VGND.n419 VGND.n369 0.123294
R1168 VGND.n325 VGND.n261 0.123268
R1169 VGND.n417 VGND.n371 0.123268
R1170 VGND.n323 VGND.n263 0.123241
R1171 VGND.n415 VGND.n373 0.123241
R1172 VGND.n321 VGND.n265 0.123213
R1173 VGND.n319 VGND.n267 0.123185
R1174 VGND.n472 VGND.n49 0.123185
R1175 VGND.n407 VGND.n382 0.123127
R1176 VGND.n322 VGND.n264 0.122488
R1177 VGND.n414 VGND.n374 0.122488
R1178 VGND.n320 VGND.n266 0.122451
R1179 VGND.n406 VGND.n383 0.122335
R1180 VGND.n404 VGND.n385 0.122295
R1181 VGND.n402 VGND.n387 0.122253
R1182 VGND.n317 VGND.n269 0.121642
R1183 VGND.n409 VGND.n380 0.121642
R1184 VGND.n349 VGND.n348 0.120386
R1185 VGND.n105 VGND.n104 0.120292
R1186 VGND.n105 VGND.n99 0.120292
R1187 VGND.n109 VGND.n99 0.120292
R1188 VGND.n110 VGND.n109 0.120292
R1189 VGND.n111 VGND.n110 0.120292
R1190 VGND.n111 VGND.n96 0.120292
R1191 VGND.n115 VGND.n96 0.120292
R1192 VGND.n116 VGND.n115 0.120292
R1193 VGND.n117 VGND.n116 0.120292
R1194 VGND.n117 VGND.n94 0.120292
R1195 VGND.n121 VGND.n94 0.120292
R1196 VGND.n122 VGND.n121 0.120292
R1197 VGND.n122 VGND.n91 0.120292
R1198 VGND.n126 VGND.n91 0.120292
R1199 VGND.n127 VGND.n126 0.120292
R1200 VGND.n128 VGND.n127 0.120292
R1201 VGND.n138 VGND.n137 0.120292
R1202 VGND.n139 VGND.n138 0.120292
R1203 VGND.n139 VGND.n86 0.120292
R1204 VGND.n143 VGND.n86 0.120292
R1205 VGND.n144 VGND.n143 0.120292
R1206 VGND.n145 VGND.n144 0.120292
R1207 VGND.n145 VGND.n83 0.120292
R1208 VGND.n149 VGND.n83 0.120292
R1209 VGND.n150 VGND.n149 0.120292
R1210 VGND.n151 VGND.n150 0.120292
R1211 VGND.n151 VGND.n81 0.120292
R1212 VGND.n155 VGND.n81 0.120292
R1213 VGND.n156 VGND.n155 0.120292
R1214 VGND.n156 VGND.n78 0.120292
R1215 VGND.n160 VGND.n78 0.120292
R1216 VGND.n161 VGND.n160 0.120292
R1217 VGND.n162 VGND.n161 0.120292
R1218 VGND.n172 VGND.n171 0.120292
R1219 VGND.n173 VGND.n172 0.120292
R1220 VGND.n173 VGND.n73 0.120292
R1221 VGND.n177 VGND.n73 0.120292
R1222 VGND.n178 VGND.n177 0.120292
R1223 VGND.n179 VGND.n178 0.120292
R1224 VGND.n179 VGND.n70 0.120292
R1225 VGND.n183 VGND.n70 0.120292
R1226 VGND.n184 VGND.n183 0.120292
R1227 VGND.n185 VGND.n184 0.120292
R1228 VGND.n185 VGND.n68 0.120292
R1229 VGND.n191 VGND.n68 0.120292
R1230 VGND.n192 VGND.n191 0.120292
R1231 VGND.n193 VGND.n192 0.120292
R1232 VGND.n193 VGND.n66 0.120292
R1233 VGND.n395 VGND.n225 0.115369
R1234 VGND.n348 VGND.n347 0.112306
R1235 VGND.n397 VGND.n396 0.111879
R1236 VGND.n396 VGND.n395 0.111186
R1237 VGND.n347 VGND.n346 0.109795
R1238 VGND.n399 VGND.n398 0.108943
R1239 VGND.n43 VGND.n42 0.108833
R1240 VGND.n398 VGND.n397 0.107764
R1241 VGND.n346 VGND.n345 0.107742
R1242 VGND.n400 VGND.n399 0.107535
R1243 VGND.n312 VGND.n270 0.107341
R1244 VGND.n401 VGND.n400 0.106725
R1245 VGND.n463 VGND.n462 0.106074
R1246 VGND.n464 VGND.n463 0.105969
R1247 VGND.n403 VGND.n402 0.1059
R1248 VGND.n465 VGND.n464 0.105163
R1249 VGND.n402 VGND.n401 0.104834
R1250 VGND.n404 VGND.n403 0.104121
R1251 VGND.n405 VGND.n404 0.103867
R1252 VGND.n466 VGND.n465 0.10332
R1253 VGND.n467 VGND.n466 0.10304
R1254 VGND.n29 VGND.n28 0.102984
R1255 VGND.n469 VGND.n468 0.102502
R1256 VGND.n408 VGND.n407 0.102274
R1257 VGND.n406 VGND.n405 0.10217
R1258 VGND.n407 VGND.n406 0.101442
R1259 VGND.n468 VGND.n467 0.101279
R1260 VGND.n318 VGND.n317 0.1005
R1261 VGND.n471 VGND.n470 0.100144
R1262 VGND.n319 VGND.n318 0.0994435
R1263 VGND.n472 VGND.n471 0.099433
R1264 VGND.n470 VGND.n469 0.0992982
R1265 VGND.n317 VGND.n316 0.0991552
R1266 VGND.n409 VGND.n408 0.0991552
R1267 VGND.n137 VGND 0.0981562
R1268 VGND.n171 VGND 0.0981562
R1269 VGND.n379 VGND.n376 0.0981562
R1270 VGND.n321 VGND.n320 0.0977932
R1271 VGND.n413 VGND.n412 0.0977932
R1272 VGND.n474 VGND.n473 0.0976284
R1273 VGND.n322 VGND.n321 0.0968228
R1274 VGND.n414 VGND.n413 0.0968228
R1275 VGND.n320 VGND.n319 0.0966929
R1276 VGND.n475 VGND.n474 0.0965648
R1277 VGND.n473 VGND.n472 0.0962384
R1278 VGND.n323 VGND.n322 0.0962186
R1279 VGND.n415 VGND.n414 0.0962186
R1280 VGND.n392 VGND.n391 0.0959861
R1281 VGND.n324 VGND.n323 0.0956231
R1282 VGND.n416 VGND.n415 0.0956231
R1283 VGND.n476 VGND.n475 0.0955348
R1284 VGND.n477 VGND.n476 0.0948777
R1285 VGND.n393 VGND.n392 0.0946781
R1286 VGND.n31 VGND.n30 0.0945657
R1287 VGND.n28 VGND.n27 0.0938949
R1288 VGND.n344 VGND.n343 0.0937672
R1289 VGND.n30 VGND.n29 0.0931452
R1290 VGND.n342 VGND.n341 0.0930016
R1291 VGND.n132 VGND 0.0929479
R1292 VGND.n166 VGND 0.0929479
R1293 VGND.n413 VGND.n375 0.0927256
R1294 VGND.n325 VGND.n324 0.0927181
R1295 VGND.n417 VGND.n416 0.0927181
R1296 VGND.n345 VGND.n344 0.0923627
R1297 VGND.n7 VGND.n5 0.0921667
R1298 VGND.n326 VGND.n325 0.0920855
R1299 VGND.n418 VGND.n417 0.0920855
R1300 VGND.n478 VGND.n477 0.0919467
R1301 VGND.n343 VGND.n342 0.0914722
R1302 VGND.n478 VGND.n44 0.0912494
R1303 VGND.n327 VGND.n326 0.091171
R1304 VGND.n419 VGND.n418 0.091171
R1305 VGND.n32 VGND.n31 0.0904148
R1306 VGND.n390 VGND.n389 0.090027
R1307 VGND.n391 VGND.n390 0.090027
R1308 VGND.n328 VGND.n327 0.0898264
R1309 VGND.n420 VGND.n419 0.0898264
R1310 VGND.n330 VGND.n329 0.0891127
R1311 VGND.n422 VGND.n421 0.0891127
R1312 VGND.n38 VGND.n37 0.0881565
R1313 VGND.n42 VGND.n41 0.0881488
R1314 VGND.n41 VGND.n40 0.0879493
R1315 VGND.n331 VGND.n330 0.0878131
R1316 VGND.n423 VGND.n422 0.0878131
R1317 VGND.n329 VGND.n328 0.0876124
R1318 VGND.n421 VGND.n420 0.0876124
R1319 VGND.n33 VGND.n32 0.0875536
R1320 VGND.n389 VGND.n388 0.0871667
R1321 VGND.n37 VGND.n36 0.0868953
R1322 VGND.n460 VGND.n59 0.0866486
R1323 VGND.n36 VGND.n35 0.0863769
R1324 VGND.n340 VGND.n339 0.0859735
R1325 VGND.n35 VGND.n34 0.0856762
R1326 VGND.n44 VGND.n5 0.085541
R1327 VGND.n388 VGND.n387 0.0855
R1328 VGND.n34 VGND.n33 0.0852048
R1329 VGND.n341 VGND.n340 0.0851591
R1330 VGND.n40 VGND.n39 0.0850588
R1331 VGND.n59 VGND.n58 0.0838333
R1332 VGND.n339 VGND.n338 0.0835966
R1333 VGND.n430 VGND.n429 0.0835966
R1334 VGND.n426 VGND.n425 0.0833636
R1335 VGND.n332 VGND.n331 0.0833488
R1336 VGND.n424 VGND.n423 0.0833488
R1337 VGND.n39 VGND.n38 0.0833488
R1338 VGND.n427 VGND.n426 0.0825455
R1339 VGND.n58 VGND.n57 0.0821667
R1340 VGND.n334 VGND.n333 0.081981
R1341 VGND.n337 VGND.n336 0.0819394
R1342 VGND.n428 VGND.n427 0.0819394
R1343 VGND.n333 VGND.n332 0.0816782
R1344 VGND.n425 VGND.n424 0.0816782
R1345 VGND.n387 VGND.n386 0.0816688
R1346 VGND.n338 VGND.n337 0.0813424
R1347 VGND.n429 VGND.n428 0.0813424
R1348 VGND.n386 VGND.n385 0.0810921
R1349 VGND.n410 VGND.n379 0.0797137
R1350 VGND.n447 VGND.n225 0.0796453
R1351 VGND.n394 VGND.n393 0.0796157
R1352 VGND.n57 VGND.n56 0.0784221
R1353 VGND.n56 VGND.n55 0.0778026
R1354 VGND.n385 VGND.n384 0.0774231
R1355 VGND.n384 VGND.n383 0.0767987
R1356 VGND.n395 VGND.n394 0.0762042
R1357 VGND.n103 VGND 0.0758148
R1358 VGND.n55 VGND.n54 0.074218
R1359 VGND.n54 VGND.n53 0.073552
R1360 VGND.n383 VGND.n382 0.0732848
R1361 VGND.n431 VGND.n357 0.0732142
R1362 VGND.n431 VGND.n430 0.0719286
R1363 VGND.n382 VGND.n381 0.0717025
R1364 VGND.n270 VGND.n269 0.0701203
R1365 VGND.n381 VGND.n380 0.0701203
R1366 VGND.n53 VGND.n52 0.0701203
R1367 VGND.n52 VGND.n51 0.068538
R1368 VGND.n51 VGND.n50 0.0669557
R1369 VGND.n269 VGND.n268 0.066858
R1370 VGND.n380 VGND.n379 0.066858
R1371 VGND.n375 VGND.n374 0.0667809
R1372 VGND.n268 VGND.n267 0.066125
R1373 VGND.n267 VGND.n266 0.0637716
R1374 VGND.n50 VGND.n49 0.0637716
R1375 VGND.n49 VGND.n48 0.063
R1376 VGND.n266 VGND.n265 0.0614756
R1377 VGND.n336 VGND.n335 0.0609482
R1378 VGND.n48 VGND.n47 0.0606852
R1379 VGND.n128 VGND 0.0603958
R1380 VGND.n131 VGND 0.0603958
R1381 VGND VGND.n132 0.0603958
R1382 VGND.n133 VGND 0.0603958
R1383 VGND.n162 VGND 0.0603958
R1384 VGND.n165 VGND 0.0603958
R1385 VGND VGND.n166 0.0603958
R1386 VGND.n167 VGND 0.0603958
R1387 VGND.n265 VGND.n264 0.0599512
R1388 VGND.n47 VGND.n46 0.0584268
R1389 VGND.n264 VGND.n263 0.0577289
R1390 VGND.n374 VGND.n373 0.0577289
R1391 VGND.n46 VGND.n45 0.0569024
R1392 VGND.n263 VGND.n262 0.0562229
R1393 VGND.n373 VGND.n372 0.0562229
R1394 VGND.n432 VGND 0.0560556
R1395 VGND.n252 VGND 0.0560556
R1396 VGND.n310 VGND 0.0560556
R1397 VGND.n292 VGND 0.0560556
R1398 VGND.n314 VGND 0.0560556
R1399 VGND.n301 VGND 0.0560556
R1400 VGND.n378 VGND 0.0560556
R1401 VGND.n446 VGND 0.0560556
R1402 VGND.n450 VGND 0.0560556
R1403 VGND.n221 VGND 0.0560556
R1404 VGND.n448 VGND.n447 0.0554302
R1405 VGND.n262 VGND.n261 0.0547169
R1406 VGND.n372 VGND.n371 0.0547169
R1407 VGND.n45 VGND.n6 0.0547169
R1408 VGND.n479 VGND.n6 0.0532108
R1409 VGND.n261 VGND.n260 0.0525833
R1410 VGND.n371 VGND.n370 0.0525833
R1411 VGND.n394 VGND.n224 0.0514752
R1412 VGND.n260 VGND.n259 0.0510952
R1413 VGND.n370 VGND.n369 0.0510952
R1414 VGND.n259 VGND.n258 0.0490294
R1415 VGND.n369 VGND.n368 0.0490294
R1416 VGND.n358 VGND.n357 0.0488306
R1417 VGND.n8 VGND.n7 0.046631
R1418 VGND.n412 VGND.n376 0.0461288
R1419 VGND.n258 VGND.n257 0.0460882
R1420 VGND.n368 VGND.n367 0.0460882
R1421 VGND.n9 VGND.n8 0.0460882
R1422 VGND.n257 VGND.n256 0.0455581
R1423 VGND.n367 VGND.n366 0.0455581
R1424 VGND.n10 VGND.n9 0.0446176
R1425 VGND.n256 VGND.n255 0.0441047
R1426 VGND.n366 VGND.n365 0.0441047
R1427 VGND.n255 VGND.n254 0.0411977
R1428 VGND.n254 VGND.n253 0.0411977
R1429 VGND.n364 VGND.n363 0.0411977
R1430 VGND.n365 VGND.n364 0.0411977
R1431 VGND.n12 VGND.n11 0.0411977
R1432 VGND.n11 VGND.n10 0.0411977
R1433 VGND.n461 VGND.n460 0.0401474
R1434 VGND.n13 VGND.n12 0.0382907
R1435 VGND.n225 VGND.n224 0.0381773
R1436 VGND.n253 VGND.n251 0.0378563
R1437 VGND.n363 VGND.n362 0.0378563
R1438 VGND.n14 VGND.n13 0.0368372
R1439 VGND.n251 VGND.n250 0.0364195
R1440 VGND.n362 VGND.n361 0.0364195
R1441 VGND.n479 VGND.n5 0.0353361
R1442 VGND.n316 VGND.n315 0.0353101
R1443 VGND.n15 VGND.n14 0.0349828
R1444 VGND.n250 VGND.n249 0.0345909
R1445 VGND.n361 VGND.n360 0.0345909
R1446 VGND.n16 VGND.n15 0.033546
R1447 VGND.n249 VGND.n248 0.0331705
R1448 VGND.n360 VGND.n359 0.0331705
R1449 VGND.n248 VGND.n247 0.03175
R1450 VGND.n359 VGND.n358 0.03175
R1451 VGND.n17 VGND.n16 0.03175
R1452 VGND.n376 VGND.n375 0.0315583
R1453 VGND.n247 VGND.n246 0.0303295
R1454 VGND.n18 VGND.n17 0.0303295
R1455 VGND.n19 VGND.n18 0.0289091
R1456 VGND.n246 VGND.n245 0.0285899
R1457 VGND VGND.n131 0.0278438
R1458 VGND VGND.n165 0.0278438
R1459 VGND.n245 VGND.n244 0.0260682
R1460 VGND.n20 VGND.n19 0.0260682
R1461 VGND.n244 VGND.n243 0.0257809
R1462 VGND.n21 VGND.n20 0.0257809
R1463 VGND.n22 VGND.n21 0.0232273
R1464 VGND.n242 VGND.n241 0.0229719
R1465 VGND.n23 VGND.n22 0.0229719
R1466 VGND.n243 VGND.n242 0.0227222
R1467 VGND.n133 VGND 0.0226354
R1468 VGND.n167 VGND 0.0226354
R1469 VGND.n241 VGND.n240 0.0201629
R1470 VGND.n25 VGND.n23 0.0199444
R1471 VGND.n240 VGND.n239 0.0185556
R1472 VGND.n239 VGND.n238 0.0171667
R1473 VGND.n223 VGND.n222 0.0169225
R1474 VGND.n412 VGND.n411 0.0158374
R1475 VGND.n238 VGND.n237 0.0157778
R1476 VGND.n237 VGND.n236 0.013
R1477 VGND.n236 VGND.n235 0.013
R1478 VGND.n235 VGND.n234 0.0102222
R1479 VGND.n26 VGND.n25 0.00911038
R1480 VGND.n234 VGND.n233 0.00874176
R1481 VGND.n356 VGND.n355 0.00816087
R1482 VGND.n355 VGND.n233 0.00744444
R1483 VGND.n335 VGND.n334 0.00285443
R1484 uo_out[0] uo_out[0].t1 984.356
R1485 uo_out[0].n0 uo_out[0].t2 582.378
R1486 uo_out[0].n1 uo_out[0].t3 566.953
R1487 uo_out[0].n8 uo_out[0].t0 478.87
R1488 uo_out[0].n1 uo_out[0].n0 424.161
R1489 uo_out[0].n3 uo_out[0].t4 294.557
R1490 uo_out[0].n3 uo_out[0].t5 211.01
R1491 uo_out[0].n2 uo_out[0].n0 204.481
R1492 uo_out[0] uo_out[0].n1 201.921
R1493 uo_out[0].n4 uo_out[0].n3 152
R1494 uo_out[0].n7 uo_out[0].n6 18.3079
R1495 uo_out[0].n5 uo_out[0].n4 17.6405
R1496 uo_out[0].n2 uo_out[0] 10.2405
R1497 uo_out[0] uo_out[0].n8 10.2405
R1498 uo_out[0].n8 uo_out[0].n7 7.5409
R1499 uo_out[0].n6 uo_out[0].n5 6.83545
R1500 uo_out[0].n7 uo_out[0].n2 5.01603
R1501 uo_out[0].n4 uo_out[0] 2.01193
R1502 uo_out[0].n6 uo_out[0] 1.0063
R1503 uo_out[0].n5 uo_out[0] 0.0793043
R1504 uo_out[1].n2 uo_out[1].t1 313.104
R1505 uo_out[1].n0 uo_out[1].t2 294.557
R1506 uo_out[1].t0 uo_out[1].n2 265.769
R1507 uo_out[1] uo_out[1].t0 262.318
R1508 uo_out[1].n0 uo_out[1].t3 211.01
R1509 uo_out[1].n1 uo_out[1].n0 152
R1510 uo_out[1].n4 uo_out[1].n1 11.6411
R1511 uo_out[1].n4 uo_out[1].n3 9.3005
R1512 uo_out[1] uo_out[1].n5 9.25399
R1513 uo_out[1].n3 uo_out[1] 7.17626
R1514 uo_out[1].n3 uo_out[1].n2 4.84898
R1515 uo_out[1].n5 uo_out[1].n4 4.5029
R1516 uo_out[1].n1 uo_out[1] 1.37896
R1517 uo_out[1].n5 uo_out[1] 0.0730806
R1518 uo_out[3].n0 uo_out[3].t1 313.104
R1519 uo_out[3].t0 uo_out[3].n0 265.769
R1520 uo_out[3] uo_out[3].t0 262.318
R1521 uo_out[3].n2 uo_out[3] 15.2115
R1522 uo_out[3].n2 uo_out[3].n1 13.8005
R1523 uo_out[3].n1 uo_out[3].n0 7.17626
R1524 uo_out[3].n1 uo_out[3] 4.84898
R1525 uo_out[3] uo_out[3].n2 0.0529194
C0 uo_out[0] VGND 9.109031f
C1 VPWR VGND 0.156964p
C2 ring_0/skullfet_inverter_16.A VGND 4.53396f
C3 ring_0/skullfet_inverter_17.A VGND 4.70918f
C4 ring_0/skullfet_inverter_15.A VGND 4.82841f
C5 ring_0/skullfet_inverter_18.A VGND 4.90629f
C6 ring_0/skullfet_inverter_14.A VGND 4.98419f
C7 ring_0/skullfet_inverter_19.A VGND 4.923029f
C8 ring_0/skullfet_inverter_13.A VGND 4.78946f
C9 ring_0/skullfet_inverter_20.A VGND 4.72064f
C10 ring_0/skullfet_inverter_12.A VGND 5.60339f
C11 ring_0/skullfet_inverter_20.Y VGND 5.35745f
C12 ring_0/skullfet_inverter_11.A VGND 4.97718f
C13 ring_0/skullfet_inverter_1.A VGND 5.16765f
C14 ring_0/skullfet_inverter_10.A VGND 5.58737f
C15 ring_0/skullfet_inverter_2.A VGND 5.65285f
C16 ring_0/skullfet_inverter_9.A VGND 4.78733f
C17 ring_0/skullfet_inverter_3.A VGND 4.92041f
C18 ring_0/skullfet_inverter_4.A VGND 4.93544f
C19 ring_0/skullfet_inverter_8.A VGND 4.94116f
C20 ring_0/skullfet_inverter_7.A VGND 4.81796f
C21 ring_0/skullfet_inverter_6.A VGND 4.53217f
C22 freq_divider_0.sky130_fd_sc_hd__tap_2_2.VPB VGND 5.57694f
.ends

