magic
tech sky130A
timestamp 1713168785
<< metal4 >>
rect 2340 -1300 4420 -1040
rect 2080 -1560 4420 -1300
rect 1560 -2080 4940 -1560
rect 1300 -3120 5200 -2080
rect 1300 -3380 2080 -3120
rect 4420 -3380 5200 -3120
rect 2860 -3900 3640 -3120
rect 1300 -3640 1820 -3380
rect 4680 -3640 5200 -3380
rect 1560 -4420 1820 -3640
rect 2600 -4160 3900 -3900
rect 4680 -4160 4940 -3640
rect 1820 -4420 2080 -3900
rect 2340 -5200 2860 -4160
rect 2080 -4680 2340 -4160
rect 2860 -4420 3120 -4160
rect 4420 -4680 4680 -3900
rect 3380 -4420 4420 -4160
rect 3640 -4680 4420 -4420
rect 2860 -5200 4160 -4680
rect 2340 -5460 2600 -5200
rect 2860 -5460 3120 -5200
rect 3380 -5460 3640 -5200
rect 3900 -5460 4160 -5200
rect 780 -8840 1040 -8580
rect 520 -8580 1300 -8320
rect 520 -8320 1560 -8060
rect 520 -8060 2080 -7800
rect 780 -7800 2600 -7540
rect 2080 -7540 3120 -7280
rect 3380 -7540 4420 -7280
rect 3900 -7800 5980 -7540
rect 4420 -8060 5980 -7800
rect 4940 -8320 5980 -8060
rect 5200 -8580 5980 -8320
rect 5460 -8840 5720 -8580
rect 2600 -7280 3900 -6760
rect 2080 -6760 3120 -6500
rect 3380 -6760 4420 -6500
rect 1560 -6500 2600 -6240
rect 3900 -6500 4940 -6240
rect 780 -6240 2340 -5980
rect 4160 -6240 5720 -5980
rect 520 -5980 1820 -5460
rect 4680 -5980 5980 -5460
rect 780 -5460 1560 -5200
rect 4940 -5460 5720 -5200
<< metal3 >>
rect 2340 -1300 4420 -1040
rect 2080 -1560 4420 -1300
rect 1560 -2080 4940 -1560
rect 1300 -3120 5200 -2080
rect 1300 -3380 2080 -3120
rect 4420 -3380 5200 -3120
rect 2860 -3900 3640 -3120
rect 1300 -3640 1820 -3380
rect 4680 -3640 5200 -3380
rect 1560 -4420 1820 -3640
rect 2600 -4160 3900 -3900
rect 4680 -4160 4940 -3640
rect 1820 -4420 2080 -3900
rect 2340 -5200 2860 -4160
rect 2080 -4680 2340 -4160
rect 2860 -4420 3120 -4160
rect 4420 -4680 4680 -3900
rect 3380 -4420 4420 -4160
rect 3640 -4680 4420 -4420
rect 2860 -5200 4160 -4680
rect 2340 -5460 2600 -5200
rect 2860 -5460 3120 -5200
rect 3380 -5460 3640 -5200
rect 3900 -5460 4160 -5200
rect 780 -8840 1040 -8580
rect 520 -8580 1300 -8320
rect 520 -8320 1560 -8060
rect 520 -8060 2080 -7800
rect 780 -7800 2600 -7540
rect 2080 -7540 3120 -7280
rect 3380 -7540 4420 -7280
rect 3900 -7800 5980 -7540
rect 4420 -8060 5980 -7800
rect 4940 -8320 5980 -8060
rect 5200 -8580 5980 -8320
rect 5460 -8840 5720 -8580
rect 2600 -7280 3900 -6760
rect 2080 -6760 3120 -6500
rect 3380 -6760 4420 -6500
rect 1560 -6500 2600 -6240
rect 3900 -6500 4940 -6240
rect 780 -6240 2340 -5980
rect 4160 -6240 5720 -5980
rect 520 -5980 1820 -5460
rect 4680 -5980 5980 -5460
rect 780 -5460 1560 -5200
rect 4940 -5460 5720 -5200
<< metal2 >>
rect 2340 -1300 4420 -1040
rect 2080 -1560 4420 -1300
rect 1560 -2080 4940 -1560
rect 1300 -3120 5200 -2080
rect 1300 -3380 2080 -3120
rect 4420 -3380 5200 -3120
rect 2860 -3900 3640 -3120
rect 1300 -3640 1820 -3380
rect 4680 -3640 5200 -3380
rect 1560 -4420 1820 -3640
rect 2600 -4160 3900 -3900
rect 4680 -4160 4940 -3640
rect 1820 -4420 2080 -3900
rect 2340 -5200 2860 -4160
rect 2080 -4680 2340 -4160
rect 2860 -4420 3120 -4160
rect 4420 -4680 4680 -3900
rect 3380 -4420 4420 -4160
rect 3640 -4680 4420 -4420
rect 2860 -5200 4160 -4680
rect 2340 -5460 2600 -5200
rect 2860 -5460 3120 -5200
rect 3380 -5460 3640 -5200
rect 3900 -5460 4160 -5200
rect 780 -8840 1040 -8580
rect 520 -8580 1300 -8320
rect 520 -8320 1560 -8060
rect 520 -8060 2080 -7800
rect 780 -7800 2600 -7540
rect 2080 -7540 3120 -7280
rect 3380 -7540 4420 -7280
rect 3900 -7800 5980 -7540
rect 4420 -8060 5980 -7800
rect 4940 -8320 5980 -8060
rect 5200 -8580 5980 -8320
rect 5460 -8840 5720 -8580
rect 2600 -7280 3900 -6760
rect 2080 -6760 3120 -6500
rect 3380 -6760 4420 -6500
rect 1560 -6500 2600 -6240
rect 3900 -6500 4940 -6240
rect 780 -6240 2340 -5980
rect 4160 -6240 5720 -5980
rect 520 -5980 1820 -5460
rect 4680 -5980 5980 -5460
rect 780 -5460 1560 -5200
rect 4940 -5460 5720 -5200
<< metal1 >>
rect 2340 -1300 4420 -1040
rect 2080 -1560 4420 -1300
rect 1560 -2080 4940 -1560
rect 1300 -3120 5200 -2080
rect 1300 -3380 2080 -3120
rect 4420 -3380 5200 -3120
rect 2860 -3900 3640 -3120
rect 1300 -3640 1820 -3380
rect 4680 -3640 5200 -3380
rect 1560 -4420 1820 -3640
rect 2600 -4160 3900 -3900
rect 4680 -4160 4940 -3640
rect 1820 -4420 2080 -3900
rect 2340 -5200 2860 -4160
rect 2080 -4680 2340 -4160
rect 2860 -4420 3120 -4160
rect 4420 -4680 4680 -3900
rect 3380 -4420 4420 -4160
rect 3640 -4680 4420 -4420
rect 2860 -5200 4160 -4680
rect 2340 -5460 2600 -5200
rect 2860 -5460 3120 -5200
rect 3380 -5460 3640 -5200
rect 3900 -5460 4160 -5200
rect 780 -8840 1040 -8580
rect 520 -8580 1300 -8320
rect 520 -8320 1560 -8060
rect 520 -8060 2080 -7800
rect 780 -7800 2600 -7540
rect 2080 -7540 3120 -7280
rect 3380 -7540 4420 -7280
rect 3900 -7800 5980 -7540
rect 4420 -8060 5980 -7800
rect 4940 -8320 5980 -8060
rect 5200 -8580 5980 -8320
rect 5460 -8840 5720 -8580
rect 2600 -7280 3900 -6760
rect 2080 -6760 3120 -6500
rect 3380 -6760 4420 -6500
rect 1560 -6500 2600 -6240
rect 3900 -6500 4940 -6240
rect 780 -6240 2340 -5980
rect 4160 -6240 5720 -5980
rect 520 -5980 1820 -5460
rect 4680 -5980 5980 -5460
rect 780 -5460 1560 -5200
rect 4940 -5460 5720 -5200
<< fillblock >>
rect 2340 -1300 4420 -1040
rect 2080 -1560 4420 -1300
rect 1560 -2080 4940 -1560
rect 1300 -3120 5200 -2080
rect 1300 -3380 2080 -3120
rect 4420 -3380 5200 -3120
rect 2860 -3900 3640 -3120
rect 1300 -3640 1820 -3380
rect 4680 -3640 5200 -3380
rect 1560 -4420 1820 -3640
rect 2600 -4160 3900 -3900
rect 4680 -4160 4940 -3640
rect 1820 -4420 2080 -3900
rect 2340 -5200 2860 -4160
rect 2080 -4680 2340 -4160
rect 2860 -4420 3120 -4160
rect 4420 -4680 4680 -3900
rect 3380 -4420 4420 -4160
rect 3640 -4680 4420 -4420
rect 2860 -5200 4160 -4680
rect 2340 -5460 2600 -5200
rect 2860 -5460 3120 -5200
rect 3380 -5460 3640 -5200
rect 3900 -5460 4160 -5200
rect 780 -8840 1040 -8580
rect 520 -8580 1300 -8320
rect 520 -8320 1560 -8060
rect 520 -8060 2080 -7800
rect 780 -7800 2600 -7540
rect 2080 -7540 3120 -7280
rect 3380 -7540 4420 -7280
rect 3900 -7800 5980 -7540
rect 4420 -8060 5980 -7800
rect 4940 -8320 5980 -8060
rect 5200 -8580 5980 -8320
rect 5460 -8840 5720 -8580
rect 2600 -7280 3900 -6760
rect 2080 -6760 3120 -6500
rect 3380 -6760 4420 -6500
rect 1560 -6500 2600 -6240
rect 3900 -6500 4940 -6240
rect 780 -6240 2340 -5980
rect 4160 -6240 5720 -5980
rect 520 -5980 1820 -5460
rect 4680 -5980 5980 -5460
rect 780 -5460 1560 -5200
rect 4940 -5460 5720 -5200
<< end >>
