magic
tech sky130A
magscale 1 2
timestamp 1712833030
<< metal1 >>
rect 18107 44260 18416 44269
rect 18107 44180 18320 44260
rect 18404 44180 18416 44260
rect 18107 44173 18416 44180
rect 12286 43628 12304 43724
rect 12400 43628 12652 43724
rect 18070 34942 18080 35018
rect 18148 34942 18158 35018
<< via1 >>
rect 18320 44180 18404 44260
rect 12304 43628 12400 43724
rect 18080 34942 18148 35018
<< metal2 >>
rect 15518 44564 15578 44574
rect 12866 44504 15518 44554
rect 12866 44502 15578 44504
rect 12866 43760 12918 44502
rect 15518 44494 15578 44502
rect 16248 44464 16312 44474
rect 14808 44400 16248 44450
rect 16986 44464 17050 44474
rect 14808 44398 16312 44400
rect 14808 43752 14860 44398
rect 16248 44390 16312 44398
rect 16736 44456 16788 44458
rect 16736 44404 16986 44456
rect 16736 43772 16788 44404
rect 16986 44390 17050 44400
rect 18320 44260 18404 44270
rect 18320 44170 18404 44180
rect 18080 43980 18140 43990
rect 18080 43890 18140 43900
rect 12282 43724 12420 43746
rect 12282 43628 12304 43724
rect 12400 43628 12420 43724
rect 12282 43606 12420 43628
rect 18080 35018 18148 35028
rect 18080 34932 18148 34942
rect 1568 22826 1788 22836
rect 1568 22546 1788 22556
rect 25650 21524 25866 21534
rect 25650 21282 25866 21292
<< via2 >>
rect 15518 44504 15578 44564
rect 16248 44400 16312 44464
rect 16986 44400 17050 44464
rect 18320 44180 18404 44260
rect 18080 43900 18140 43980
rect 12304 43628 12400 43724
rect 18082 34946 18142 35016
rect 1568 22556 1788 22826
rect 25650 21292 25866 21524
<< metal3 >>
rect 15492 44568 15602 44582
rect 15492 44504 15518 44568
rect 15582 44504 15602 44568
rect 15492 44484 15602 44504
rect 16226 44464 16336 44480
rect 16226 44400 16248 44464
rect 16312 44400 16336 44464
rect 16226 44382 16336 44400
rect 16968 44464 17078 44482
rect 16968 44400 16986 44464
rect 17050 44400 17078 44464
rect 16968 44384 17078 44400
rect 18306 44260 18418 44278
rect 18306 44180 18320 44260
rect 18404 44180 18418 44260
rect 18306 44162 18418 44180
rect 18060 43980 18160 44000
rect 18060 43900 18078 43980
rect 18142 43900 18160 43980
rect 18060 43880 18160 43900
rect 12282 43729 12420 43746
rect 12282 43623 12299 43729
rect 12405 43623 12420 43729
rect 12282 43606 12420 43623
rect 18054 34934 18064 35028
rect 18168 34934 18178 35028
rect 1558 22826 1798 22831
rect 1558 22556 1568 22826
rect 1788 22556 1798 22826
rect 1558 22551 1798 22556
rect 25640 21524 25876 21529
rect 25640 21292 25650 21524
rect 25866 21292 25876 21524
rect 25640 21287 25876 21292
<< via3 >>
rect 15518 44564 15582 44568
rect 15518 44504 15578 44564
rect 15578 44504 15582 44564
rect 16248 44400 16312 44464
rect 16986 44400 17050 44464
rect 18320 44180 18404 44260
rect 18078 43900 18080 43980
rect 18080 43900 18140 43980
rect 18140 43900 18142 43980
rect 12299 43724 12405 43729
rect 12299 43628 12304 43724
rect 12304 43628 12400 43724
rect 12400 43628 12405 43724
rect 12299 43623 12405 43628
rect 18064 35016 18168 35028
rect 18064 34946 18082 35016
rect 18082 34946 18142 35016
rect 18142 34946 18168 35016
rect 18064 34934 18168 34946
rect 1568 22556 1788 22826
rect 25650 21292 25866 21524
<< metal4 >>
rect 798 44610 858 45152
rect 1534 44610 1594 45152
rect 2270 44610 2330 45152
rect 3006 44610 3066 45152
rect 3742 44610 3802 45152
rect 4478 44610 4538 45152
rect 5214 44610 5274 45152
rect 5950 44610 6010 45152
rect 6686 44610 6746 45152
rect 7422 44610 7482 45152
rect 8158 44610 8218 45152
rect 8894 44610 8954 45152
rect 9630 44610 9690 45152
rect 10366 44610 10426 45152
rect 11102 44610 11162 45152
rect 11838 45008 11898 45152
rect 11836 44952 11898 45008
rect 11836 44610 11896 44952
rect 12574 44610 12634 45152
rect 13310 44610 13370 45152
rect 14046 44610 14106 45152
rect 14782 44610 14842 45152
rect 798 44550 14842 44610
rect 15518 44569 15578 45152
rect 15517 44568 15583 44569
rect 200 44140 500 44152
rect 798 44140 858 44550
rect 15517 44504 15518 44568
rect 15582 44504 15583 44568
rect 15517 44503 15583 44504
rect 15518 44500 15578 44503
rect 16254 44465 16314 45152
rect 16990 45080 17050 45152
rect 16990 44952 17052 45080
rect 16992 44465 17052 44952
rect 16247 44464 16314 44465
rect 16247 44400 16248 44464
rect 16312 44400 16314 44464
rect 16247 44399 16314 44400
rect 16985 44464 17052 44465
rect 16985 44400 16986 44464
rect 17050 44400 17052 44464
rect 17726 44506 17786 45152
rect 18462 44952 18522 45152
rect 19198 44952 19258 45152
rect 19934 44952 19994 45152
rect 20670 44952 20730 45152
rect 21406 44952 21466 45152
rect 22142 44952 22202 45152
rect 22878 44952 22938 45152
rect 23614 44952 23674 45152
rect 24350 44952 24410 45152
rect 25086 44952 25146 45152
rect 25822 44952 25882 45152
rect 26558 44952 26618 45152
rect 27294 44952 27354 45152
rect 28030 44952 28090 45152
rect 28766 44952 28826 45152
rect 29502 44952 29562 45152
rect 30238 44952 30298 45152
rect 30974 44952 31034 45152
rect 31710 44952 31770 45152
rect 17726 44446 18142 44506
rect 16985 44399 17052 44400
rect 16254 44396 16314 44399
rect 16992 44396 17052 44399
rect 200 44080 858 44140
rect 200 43724 500 44080
rect 18082 44000 18142 44446
rect 18307 44260 31938 44269
rect 18307 44180 18320 44260
rect 18404 44180 31938 44260
rect 18307 44173 31938 44180
rect 31768 44152 31938 44173
rect 31768 44050 32100 44152
rect 18060 43980 18160 44000
rect 18060 43900 18078 43980
rect 18142 43900 18160 43980
rect 18060 43880 18160 43900
rect 12298 43729 12406 43730
rect 12298 43724 12299 43729
rect 200 43628 12299 43724
rect 200 22862 500 43628
rect 12298 43623 12299 43628
rect 12405 43623 12406 43729
rect 12298 43622 12406 43623
rect 18082 35029 18142 43880
rect 18063 35028 18169 35029
rect 18063 34934 18064 35028
rect 18168 34934 18169 35028
rect 18063 34933 18169 34934
rect 18082 34928 18142 34933
rect 200 22826 1810 22862
rect 200 22556 1568 22826
rect 1788 22556 1810 22826
rect 200 22538 1810 22556
rect 200 1000 500 22538
rect 31800 21540 32100 44050
rect 25642 21524 32100 21540
rect 25642 21292 25650 21524
rect 25866 21292 32100 21524
rect 25642 21260 32100 21292
rect 31800 1000 32100 21260
use freq_divider  freq_divider_0
timestamp 1712832449
transform -1 0 22072 0 1 43628
box 3864 0 9552 640
use ring  ring_0
timestamp 1712778044
transform 1 0 16088 0 1 22922
box -14600 -14600 14600 14600
<< labels >>
flabel metal4 s 5950 44952 6010 45152 0 FreeSans 480 90 0 0 uio_oe[0]
port 19 nsew signal output
flabel metal4 s 5214 44952 5274 45152 0 FreeSans 480 90 0 0 uio_oe[1]
port 20 nsew signal output
flabel metal4 s 4478 44952 4538 45152 0 FreeSans 480 90 0 0 uio_oe[2]
port 21 nsew signal output
flabel metal4 s 3742 44952 3802 45152 0 FreeSans 480 90 0 0 uio_oe[3]
port 22 nsew signal output
flabel metal4 s 3006 44952 3066 45152 0 FreeSans 480 90 0 0 uio_oe[4]
port 23 nsew signal output
flabel metal4 s 2270 44952 2330 45152 0 FreeSans 480 90 0 0 uio_oe[5]
port 24 nsew signal output
flabel metal4 s 1534 44952 1594 45152 0 FreeSans 480 90 0 0 uio_oe[6]
port 25 nsew signal output
flabel metal4 s 798 44952 858 45152 0 FreeSans 480 90 0 0 uio_oe[7]
port 26 nsew signal output
flabel metal4 s 11838 44952 11898 45152 0 FreeSans 480 90 0 0 uio_out[0]
port 27 nsew signal output
flabel metal4 s 11102 44952 11162 45152 0 FreeSans 480 90 0 0 uio_out[1]
port 28 nsew signal output
flabel metal4 s 10366 44952 10426 45152 0 FreeSans 480 90 0 0 uio_out[2]
port 29 nsew signal output
flabel metal4 s 9630 44952 9690 45152 0 FreeSans 480 90 0 0 uio_out[3]
port 30 nsew signal output
flabel metal4 s 8894 44952 8954 45152 0 FreeSans 480 90 0 0 uio_out[4]
port 31 nsew signal output
flabel metal4 s 8158 44952 8218 45152 0 FreeSans 480 90 0 0 uio_out[5]
port 32 nsew signal output
flabel metal4 s 7422 44952 7482 45152 0 FreeSans 480 90 0 0 uio_out[6]
port 33 nsew signal output
flabel metal4 s 6686 44952 6746 45152 0 FreeSans 480 90 0 0 uio_out[7]
port 34 nsew signal output
flabel metal4 s 14782 44952 14842 45152 0 FreeSans 480 90 0 0 uo_out[4]
port 39 nsew signal output
flabel metal4 s 14046 44952 14106 45152 0 FreeSans 480 90 0 0 uo_out[5]
port 40 nsew signal output
flabel metal4 s 13310 44952 13370 45152 0 FreeSans 480 90 0 0 uo_out[6]
port 41 nsew signal output
flabel metal4 s 12574 44952 12634 45152 0 FreeSans 480 90 0 0 uo_out[7]
port 42 nsew signal output
flabel metal4 31800 1000 32100 44152 1 FreeSans 2 0 0 0 VPWR
port 43 nsew power bidirectional
flabel metal4 200 1000 500 44152 1 FreeSans 2 0 0 0 VGND
port 44 nsew ground bidirectional
flabel metal4 s 16254 44952 16314 45152 0 FreeSans 480 90 0 0 uo_out[2]
port 37 nsew signal output
flabel metal4 s 16990 44952 17050 45152 0 FreeSans 480 90 0 0 uo_out[1]
port 36 nsew signal output
flabel metal4 s 17726 44952 17786 45152 0 FreeSans 480 90 0 0 uo_out[0]
port 35 nsew signal output
flabel metal4 s 18462 44952 18522 45152 0 FreeSans 480 90 0 0 uio_in[7]
port 18 nsew signal input
flabel metal4 s 19198 44952 19258 45152 0 FreeSans 480 90 0 0 uio_in[6]
port 17 nsew signal input
flabel metal4 s 19934 44952 19994 45152 0 FreeSans 480 90 0 0 uio_in[5]
port 16 nsew signal input
flabel metal4 s 20670 44952 20730 45152 0 FreeSans 480 90 0 0 uio_in[4]
port 15 nsew signal input
flabel metal4 s 21406 44952 21466 45152 0 FreeSans 480 90 0 0 uio_in[3]
port 14 nsew signal input
flabel metal4 s 22142 44952 22202 45152 0 FreeSans 480 90 0 0 uio_in[2]
port 13 nsew signal input
flabel metal4 s 22878 44952 22938 45152 0 FreeSans 480 90 0 0 uio_in[1]
port 12 nsew signal input
flabel metal4 s 23614 44952 23674 45152 0 FreeSans 480 90 0 0 uio_in[0]
port 11 nsew signal input
flabel metal4 s 24350 44952 24410 45152 0 FreeSans 480 90 0 0 ui_in[7]
port 10 nsew signal input
flabel metal4 s 25086 44952 25146 45152 0 FreeSans 480 90 0 0 ui_in[6]
port 9 nsew signal input
flabel metal4 s 25822 44952 25882 45152 0 FreeSans 480 90 0 0 ui_in[5]
port 8 nsew signal input
flabel metal4 s 26558 44952 26618 45152 0 FreeSans 480 90 0 0 ui_in[4]
port 7 nsew signal input
flabel metal4 s 27294 44952 27354 45152 0 FreeSans 480 90 0 0 ui_in[3]
port 6 nsew signal input
flabel metal4 s 28030 44952 28090 45152 0 FreeSans 480 90 0 0 ui_in[2]
port 5 nsew signal input
flabel metal4 s 28766 44952 28826 45152 0 FreeSans 480 90 0 0 ui_in[1]
port 4 nsew signal input
flabel metal4 s 29502 44952 29562 45152 0 FreeSans 480 90 0 0 ui_in[0]
port 3 nsew signal input
flabel metal4 s 30238 44952 30298 45152 0 FreeSans 480 90 0 0 rst_n
port 2 nsew signal input
flabel metal4 s 31710 44952 31770 45152 0 FreeSans 480 90 0 0 ena
port 1 nsew signal input
flabel metal4 s 30974 44952 31034 45152 0 FreeSans 480 90 0 0 clk
port 0 nsew signal input
flabel metal4 s 15518 44952 15578 45152 0 FreeSans 480 90 0 0 uo_out[3]
port 38 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
